 GITCRYPT Ih�C��
��k"�v��B�z ��3��ߎ@��j�d�01(k�U1� �/��0����k�k�d�#�@���l��M�,�.�����b�ƫ!P��l�{�=��o�|���=s_eMa����HԆ"�rW+ߓ
��.�Sc�^�&�7)�BM�`7�#��*��Ћ�A��O��*�^h<^W(���&��m���VV�S�ץ��6&��#�̀ƴ�:�	��&�0/�B������Y�R�s�q���z�,��}��}�Ӧ�&V���o��Ts�*���h��c�-ܢ��zg�c��<��՗�;{�S�n]�J>���� �k^���g[��z�b�Rʊ�;^(�fe��mb\���S�XT�<�EI$M.��2���n��F��15~�3A���D=���N�	M���"�̈p��n��?k*X����~�W�_t���Η�s�S����ׯ�\�#�jJ�D�g��_��$�͈�3:�D�wԏJ�N�3�/䓹��둫"܍�	o��S�c���о������t����BX���x���l�E���s���?�D�B9��ŝ�tV.��cq{��=�
DR��4�Y�7�t?ӽk2H�������;������[%W;�QG�bvxͧ���I�Z�԰CVr��?0�<f��3`�+9��Ni�|>�!诀�9�S�T	UD�Y�
� �����s����.q�dM\1�
��W��<���ahiZm��\�._'q-<t��=�D��� ������;�J_�m��P�8����]`�.��*zѴo
��T�M����ѱ���yo�nU�����MN��"�KiɆDp+ҧ��ϰ��!@�˒�����ςf���
��H��͉3BWnH���G��u��y9H$4�8�z��}"�6-sI�<6�2�d�dh�	�J���b,5�NV)�����+�S��_�&d҆c�K�{��@h'�%�r���B���йȏ^Ɏ�'���q5�u;�9琟)�U�.�pB*P�phv�',���U�	���V������q���<v.0n+���)��`CJ�:�Z�K:�v4�)��ȗ�@Թ��"�V��Ѥ�PĭY^���*?�,@�Gbc�D��d'9��hCKĖMN�C�7����Ȱ�����,���n��i�D�{�F!W�_?[��� ��i�?���um�~[�؍Se)����Ι����ծ�N�����#^���Qk<�8$Ao1Dߞ��WѾ(����j9S(�,��قÐ8�l��R[\+%���glս𤛦>�Q�N�ܢ�=��_:m�Č�ԐؐK�@4��gZ��Bx�Ͻ;H2�.�ۃ6���Ob�.~�?xF�����H�zr��gȑ�������Q�կ��x�_"�m��a��]hD����zh�b��dJ�n d���
O���(���>$(���ޟy�O�L��z�ey���ǵ�)2��u���	�����#u��3Y�H>�b���鲙��Ď�w��	)'�4�Ȝm���=�_�8�s"���b��fq�	��A�"P֖��~���㏺�p�v��D��2%=��&!�+���>�H���<;�v@iթ��S��p)�Xժ�����<���6K�#E�o�#�-���&���B@om~e�Eg����C�r��s����^f��e|�p�o���x�J�0Ɇ�?��C����?v΅�$RM�B5�G�(�V��?UP�U�ދiħ$�/y�^
ҹ����m/N�@����sP����c��(�y攡A#x�g-�T� < &Y>����KW�,Di�.�Z����sWtaS7�^��LO�2s I��*�N(h���"=Z�Nw3̵�UvȚ����m��=��]�ԌAQ+"�'�������}�����
ʹ�*K���1?�� ����ʱ� ���|ɖ�Yx��s�(u��l���+ޢ�3�zi"-$���λw�㛌�\��	Z^s"-�������CE�j������	����(�.��^Plxu���mDr�k��u���w�hb�O��!���:oN�jA8�O��= E�XI�P�N%�\�;B�ԝ�{���h���[��L��e3Y����0#\�WMd
7��%�=G ���GA�ɗ��b\S��&1d�"NB���MZK��Rԓ����aX������X��	����6{�n�!�X��fkH�ʖDd�'Ųm�D��c��������z(�sC+��g�g�<6[���@P������<rzgg�8\*�\ח��e��������������e�,&��U9�F9r hV�:+�F��ܚ�� g�K�`�}g��GS'Yb�4M��ϫ�!�M�>�u�*���y~VΔZ�	0���{T?���3���3@�	0_�,/4@�|e'�'�+�zKf�U׌�".��7+�z�yH��,��/��|�d!�oL��\��0!��U��W���队�dh���j4F�}�&bQ ���y�00�:��`�F�
"8E�6��wj��R#���%T�m8���.�:�XI���.]�X�W���r�?��,˿��vb�K��8:����m}������Z$T޺g�\�
�,�<���ry/N@G�̓�X�Sc
���՚ё���a��f8~�~�� �gՄ-�Ϧ����}N!��zP��)��wޗ���<�g`�O�vk���J?���W�{�<�;Š;�v^ꤙK�ta�{�Du�ã���.��=�PȊ���'o�"���H����~*s�̣��}�����P
�.�`�,z��.�K�yUbW�z�ʝ�|�Yk2����,��s��>@xUЬA�R��1,��z�?cl�J�wo�~��$8�V��U� ��Z��?��W�v�c���Z���r�\��@�͟��OІ�_�$K�U��m������)ͣ�m�kwo�j���r�Ԟ- ���̄�I�VHu,��(�\��;�cǌ"���;�_�2u�n<��C^�aH��,�X�
Jl`L|#�4�D�a��.�=KፏV�}�`�M�GNO}�Z}��ȲP�}T�W�t,��c'
L�?�� ��܎��=C"�Te}8�I�Kʒ���ѓ����R�-��ϴ�T�
3xl�$ �n����>Hm�e�7�>��a������z*4[{�,9/�<{z�m���ar�̆qϯb �im���*����<d��"�hw��q|�j�
i�Kx��9U� ��x��cMY� Yu�$HҨ̠������ts�*�LY���Z��@��T�y@�&�LE�:#�}P�OQ\�7h��I	E=�����,�(��.��G�sjp��
�䫗��
'����h	��]~��	+䟜�3ǚ)}���J�]�����pІ�5�>imaKx�����'���Q��[��*��������3���� mc����7���8�\��[�E`���/;(F/�B�W��h�(��O.��k���3��O(ϣ�����l�CC�.�˗�U`�b�6��SjOP����P�{;+"��q�p"%5S̪;9�n���%��@ �4��3. �_;�a�>�^�����&�4A�Ɲ���r��qh[����p��[4������?���U�30��"�)f^���V��p��.�)� �E���2
=�L�S�U�ҫ�����-<Q�v"�M:������Ġ�u��q Kr�%�#����Ven�3�(f����b��<�rJ�pa���RM����
��w g}��Nu떭�0I��Mt�l�o؊pƧ&��8���+�e8�l�vnl�Z4j+4��ޘ�QQ�{;9�*��'π=Ү�#��g�ӱ��I�Wߤv���|VUE��w�$������	��#�A!<l@o��5��/�V�G5笝�$��:P�(Z~)����,��xƊ��M��hDI�iQ+�s����aY0�x���%AA��A�����8�Ս����z�m���[~�	�J`�M� p���36:]p�n1�]C�b/�tp��K(���;�_���	0hsN"��J@"���f���{#�`�M��t*뭣�;	p����l1���pUZߕ�j�ӘX�2���P���\rK��p.O,E;NRf\�V�}�4ۼu��Zv��,���@���� �Yg=��X���s�u=��SJ�Ѥn�T��p���e���S�Yc0�;�����G6��H�Hm�.����C�x<��<�ݎ���¼���s�"���ypt�5�����~)j�m�š��1i]$㊕EjP���E΅ ��s���jIɶ��K�fv/�\��7-j3a�F& P�?�����c��渓�f��,�×�@=Oѻ�bF_3)��"�����}�,D�gԹ��w#���,����=�ʫ*ţ�Qcm%�Q�S�T�l=�E���ߧ��e��O�0<ŧ"��j�s���L\ྥC��e~.I���'�%�2k����6M�ƭ��O��.��r�{-Z�"b�,��y���D ��@�N���-�&�E'��ґk�s�̩ë�tU-]�-�����R���G��ٝd^�J������ 8l��¬�屩�xf.0���t�JsTb���VX���Է��0�(��I3��VbO��wm��pr�����*p�?&�ǿ��M���ƅYN`%I���M���-�`:n2ښ�w��bT���b>L<f��?9���o�j,�$YA�T��:�v ���(o��5�W�%sWj�N�(��O6��B��p�ބ9�:B'>E��-ً�:�̇��j��0�f(��"�,:49�Y���j��}��ؔ��K�x�s������j�d��HO�X�SH���W�S��9��X��H�d��Ǫ�"B2�"�[��83}����Bt�`�/Q,��{<*v[��*\��V5*� �x�ܥLl��@�O���@�f�F�Z|Q�1���.#^����!C�c�� ����AgE���c����r1YdV���K��y_l��8u���-�8�N@����s�r�3 �~�35��ɠ���6&3F~����|��іE�p�1��x�U%�l:kť�y5s6!U�l>��1�T�H`7�����FF�����|l=i�<a=�r��P#�W�Tґ#�NTBċ�e�Z����pW,�6�%� ���`|�,�NZ[���1�s�;�&�{��ǁ�6��k�Q������Tc�}Q}
������i���ZNh ��\pFh�]���^6�3��sv��S��9��<���!݁rv��'>��!������JX�׈��B����tq�r�hi2�{HI����eN/C��g�c�QT�v�\�2w�'f)�Q(��'g����!��n�����@\-&>���#�ͮE/P��AQ��:6BVO�O
=��k�e����t�t�� �����	�u�����6LG�>xc��_���l�g�dr���
���w0�̏[�B�(�A�j.v�K�-��1r�Z�Z닞��N�"GSgR�3	g�޲%n}x�E�%�-��><c����C�RYI�޾��,͓�ݨbo��:��ez���]TI9w�;U���QT�<�eXr8�����g�h��^��dm�ԍ���=wz�~�
�	BO�[X=���� X޴z��*�Y"?P��D���|��;���g��q�~�Ȍ>S����� �c����3��z��i	�p�BR�vZ㠠���>�eˡ��5k단en��"'w�ga��Z��iC��#�FxΎ/��3�ǵ�P�d	��ճ//�����#@B�\��JsTX��V C}�v�ٗ�:(]�#��n6T�۞o ���/�e@�������t<b�i�G��u��njl.�g�(X�����U��
:�h��#�g��� �#�n1R��1�	(��<ǣ�=�|�:����,�zS灏غHՠF�w���_-���A�a��l_�f!�}y;�n ���t�]�qf�JTpQ(O��I�t���D�w;\s�r�����vh�p\��Z���fr��`�^�`���^N�ǔ�7���R���O�Er��G��.Iwur��z2��̈́Гh��0@����Svj9-1��~c�-}�p���5N�t�1)�G0)0�Blϐ� ┼���D,J���ާ>�B$��OM%���E�+�ר�c�����K�}�����}��;O3*R��X0!M�e&�R1��	��]�]�Z_��X:��н�����k���h�l�5��l��d��&v�l���F=�ޣk���;�W��`�oٕ[;��X60��VB�k���o	�@�WG����Ԣ��������#*[��u����k�6}EQ!���5F��=��VP�q�[��#&mh���4P�N���i�0�
9������կ�c��E[>p}��X����%��~�y���� ?谭�M�F&s����o�(�����-�̞v'�p}BǤ��짰��]+��v,IjClwJV����K��u�I�r
ز\g�*����O�d����w$�U��U���v�8�Y�5�(���2��X��=��ǚ[/����6O����|��sKot�Ǡ>�[�E��Nl�`��|�
�s���_�mR�����"��x3�Q���A(���3��cJ�j�Svwf����z�<7��y'�~��hg�+ܘb~'��㔸���D���w�4=�=�k��U
�Tm%�j�n�Z�`��Y��Q�qu����o���TrkM�m�ͅ t�g��s��K���9�R�.�(�O9R=����Z���R�X1�D|V!WP�ξ��Hz�P�	 ��V�g����^��w�#Z�V�{I%�$$B��*x*=�틄��u�q�?�d;h���<��(BeFI��֋^F�/H#�'#����6!j�5��V��Q�=�*�w;�u���QV���.0l[�-tv,��v�T���uR��v��Fu�';1��q�^�_%9^��]/�{��J�`�X�F�d�A����`���*!��RQ_I��������XI��h���]�<Μ�:.Πl���'���^�G��m5γR�9'@C���f�C���$�����}-Yd6Zk�����й�����{�D�"x�'��-�ذҞ,���{�$�P @h݅� �^����'�cF���Tf�w+Գ���[y��b�K�rRp��@����x:�\�kl[,�++����K�Ӂ���_��@ѧ�NB#�,��K4��@$0<��`?wػD���j���*��ׂD��^�tk���ASp.�s�����b�(�P�~��v�Iz��_��С�<�