 GITCRYPT w���L3�ط�.��Rş���a��ݵ+�(D+�_��������%�l�Q��(�RW6�g��J_̖#�[��'B���@��cj�?ߒ9���	��ހ<²��$CJ����=[�5d8��`���������tU�҉��}WX�Q;=(�|�kO�^�h�g��F`6t�f�x^�5��?�ߔe�"�-*r�ɨ#.�R��?�]F����~-E'�A�O�PLV�/���y^G���Ɵ�x�Pg0l�2-gI����/�!2����=P��5�a���v�ňE��9���kFv�嬂�'�c,J_� �Y���M/��}��?�ݎ���TbUi��d9��Bڽ�	r������V���W�UK��?���a����,{�(��@/�T�&�o�r�A�t��g��w��ef6��_Y$���̱���z�<n��/���-J�<�Cl0�F�ub�h1��yS��ד��FF`��L7�j�1���0]�ڽ�B-N�'CP�6P�ηs�sXe�%�Tw���(��I�!a!�Oj?����3�s���mP�	fy�La�1���cl��`0^�1�7gq�$!��bAL=r���jk��o�J��@�Ky-Q�"����E����z@�΍���q�>�k�y���c5C��|�&l�a�����{mVuAH�
�L�
�S��'�J-���,|g*�ޅJ�,�SKz���	Dl-�:��C~�D���@�I�1�5�n��5&�ɖ�����j/<F��5.�7z��oV ޽x�G�7=HV���)�Q�S"�&��d�L0P�;�Y��AKѭwRF� t�*d1�� �t��'z��M9V ������xbm
�ۆ#��8�P�[��7	}�)�dM��������~�&y�������ۿ��@����R�dD#� �!����B�w6���on��z�����Q��n{��żŠ�u/�)�@�u|?�npE8���D?��&D��g��d�BGX߸)s���^4�|{K2�����>�S��0CW/�,Ũ;�S�8KO||	lA)r`����h=��/�W�C0\������F���~��h���q(Gh: ������7��
��*!�p��O�;-���Z��
*��9��R��ͫH�T�n:��Rg��Q]�G�)�ATQ�!�y�P$)4���^���J,��G�o�Xa9�nI_fd��Iq�d�X�}��� ���|1�̎�9F1��9Q�ϩ�)�����7?>���4A���;&�$$�o%3��	8��������f1A�}V�g@���l"+i��5�p!Q��q��,r�qjB꜎� :��=����&�f)|N`�2`Oi��e�'q�Y؟�MzRV&,C���n�|�=D��c��o+7<g0�?���wQ�y����ۀ� ���:�W1X s1gO'j�S'�xH�'od2*���Rf�� O�+8��y�����B�+?�`C#��y�s+~�8��n�#�޻�`�9#ݖ���Ǒ��J��%�b�dd�*��-t}i2n~�!
�#�6��tRR�f�wkJ��e�c�rx`&e�ÿ(c\c��CS: l0�g�#�VD.��q��w}���E���T-z�f����"ԡ�1�s��)h� j�L�:��?.�����V���� ����*n���K�ġ�"�oc�1}�H�g�6����.G���Lѡ&7>�0[��^_l/WAR��տ��h��҆|y�J��K���� ��s;�B���
�b�e�
3�
W=M��x����M6Dm�+����s��Qd�-�1hH�+`��FuuY�8�¸p'r��8}V�9����H��"I�l"�u��#��Q@�~T�X]i�c�����A�3yG��bJ��mNOp䑭��r����\ ���x�C��'-�3w�!I䁣�"8���)��4��>=*���(�Qd$����5��C8�;��ا�mV�BR�/�]^,)&�@�ʦ�,��� a/Q�Î8�ʚ^�O "�� R��������ﺀUO�|`ŒyxB-UN��n���"�+=Wv���ϗ`pr�5z�a�i��]�*���Б�F�NG��~ż�52*�g����}y�g��Ţ%�;I����U�Z�6��(A��2	?����-���<�ω9 J�	�'��Fhl�� o�F�J|�sA�X���K�9��i�\���ؤP~�e^k:��Y�k���+��o�&�k�L�D�[,�޹������+t�J�g�`�d]�/��0���s���������o�����:K�~�	QP��
��eVJ���kcQ���͑N�(�jc�)���3ԯ/n���c�7I�G�6�6i��k�T[8��Ss"C�5t��
�3��Q�nת�k�H��2�PDRDUr� ���S0��;�2��\���Z�Yv1��8�����N������Ѧ"<��B�ɱ�$����S��k���՝��tEE�I�ԏ|M�&����2�U��V�BDQ�͵���]Щ�$M�V:�VT6���!	�=b���?���1�����Vf����ȬS��eC�����%}m���G�:mmv�
8K����:3�Rsij�k�6~���U�����jM�O*H�#�x�$���s�Z){�M?; ����9Tҏ�SR5����b-�&��9�ER��D��p����Ѯ���}�s��Zr�G�l!,�u`
��]��C��}d˛�\|��� �`�R��
�¦�s%�QJ�@+�8�)����-��y;�`��&�0�s��F�Z[Ò��<pW,I�,S&J� ��K�_h[p�&6��:E������-s�nS�ɞ�b�d�*րl���M,�ne�f�h���f�I�X�1Z��&4`1PW�e$�!�4�)�_\���w��q�=��'������}q�R@rצ��JP~�C:�y�mk�M[�S�-�������F��-��F]���r���p�d|���d�_4�}OIA������]��$�Z���mT���E򲿶��:�(�Nh0;�i�;�Z�[w�>�w�����/L!nm�%/�ٸ�a]�PM[��ozP3#PN�S��ȗ��,�B����AR��I�e�sV����uE��J�U�d�Kp��YX#��;�n����;��-��P@�[�ዛ?�µ���,�FQ���q��!4�Э��Fm-2)�#'%Ň��6_����σ�� 9�ts��x[6�L��Y��"�}ŷz���Z�B2����yW�T�N��wT���C�iXdV'��؊)���{�0*�I9T�/P��j@ ����3f	o Z!-rŘ�`��	;r�!g�K�e36}y����KK�y�W��,:��ք�9,� 9���=]Mq`E�e�����}��":r.��$�=/l�ҍ�x���B�T!��NK	56��~Ki�M�ݳ�
b�ոNQq�&��!��~�΂��v����κ��Db���mTk�rD�ݻl��͙��[@I9 ��+�f��Ô�;me��5J��n�e
���9�(���)}0;�i4J忴*�)ڹ�+z��IN'����劅EO����
h���kb����"����?STI肢��pW��tJ�8m�a��-&^+�}o!=$|�'Uq;+�;[+|@:��S�^�N���.���Yz��� <q�s��_��t���'3�2�XK-|��0L|���S�O�t*����m������i=�Ɲn-��?T��]���h���O�#�I�(��-�)��MX�2�O���s���J�;�g*'+�����69���U�"F�b�Q}K�5j�
8B@f��I�6k%T��^��5�1L9����=�T�M5��!S�9���Wx�q���B3� ��>�=�W?�Z�Md ���0m��\0c�)ـ���	<l)�T�����$0_���<C݃F}��f8����qj��|����*`��n���66Z|+�/�C���K�p�O	^^��\q�
�RL����ߐ�w�XM~�ƴ9x�=%���Dm���2��d�@%w������j��L�d�uS��-����c�AI����˼-|4#+ �(z�C�$�(�Iڭ��<�M]����( �Ǖ�X������lx����v�VV����b���>=��3ǒB1]��r�y��͚��`�%�қ��ц�J��
�~Y���u���'�lc8�⫍`p@�Ơ��-:�?\�"�U"�T*^u%EYO)����]6��N��u���C&Q>T4p[s+-Ҹ�ަȸM��K,)����m��O��344�pb��=ߖ����oj};��Q�JR�38)~�0��2�^p��TϘ�\�N/e�A��������N�$)(kJB����ͪG�����	E�=�i�"��t|�nq����#�@/�2�������� (z�<kqyk��p�YU�Si$�S���P���׮=l�"tj�U)��д2(�+�������Ǧ=KV������#1!�z��I��=�&0K��g�����-��A����49�*4"G�a���p�%��n�Ð�����^��E89�`�aˑ �by9|d���x�\�v�7�NY�"�^m'�ʄ�F_M	>��0K��7E�b��F�k�˔�~����[)8����R��H��Z)�i}"��4�x㫊!:5�JY��uN�M���Vy�B�T���K��8��e:K���9V��e���Z�ܘ ��{�����>K�T���5�����@:8s���os�FΌ��O5U�␭0^z� �����ٖL�	�)�I��+ XKz�	���v3{3����(Q �ɇzS��� gS�ʸ�&���\|I|�էtשp@����3����d����Z �=I�Z�¢��ݲ~��H�3]���3/�[�cW���dPQo  ɭj���"�F�:e����V�e["�Q>^��'~�$uH�'�!��<�x��v�����v��~�M��\gB�s����x�
N:橂�D)76��6G��j���ފ����_����!к�T@.!��ؼv�����`H`��u\�X�l�H~K�[�[�T�V���a�0�o���a>NHBC2�E�fM=���"���Gkfo��j����&�Ft�p�rx� 6��f}��V�ϙ#K@��:��F��`�rT�����'{zTJlv��m�<ß� T�$h.��J��B���K��z�x��v�oY���d\xm�,���=� �mi_$�6${�gݜ�b��]>���hfCG�:	�$��W,�5$l�o��L��G��!�p4������� �:���2�bnB�y�g\]Դ���f.��E��A����j�����Zi5����:�X�
VV���m59�a����6h�%�d�{����@��~��A� ��(L<A�RQ��7��W{���Xb��(i�i���m@�m��9�eN	rï-�t�R��bfk��d�ֱ�cᷣ��C�4^;	�^*Օ�f�[���	�yH��7�k�Qk�Z�t͝����&��hs`3kaֹ�'�5��kE��92����������������w�-@(N�RA��S�-K-��9�s����X5J�բ����N��Md��r\�۝�RjN2+ <�ia��}�|������A��˱o7ƲX�aJ�읷`ÿ@ob���7��sg����׎|{Yu�Q H��\k�_jk`R?NM�9�������[
��X+�e�<�\�>^�|
'#U�Hh���x�{ʢD�����v�w�x×
���4oں~p �_���k�a�n������I������YB}���х֚�J��a�=l��֨�?06=��"j�3����`9xׅ������Visa!K}��T�JsZ�>_�D6�+]f���s,W\JFAP1��l8Ή��\0�aei\��V�7�AD#�@�1N�V*��^����SM &������@�*lFF�:�ʙ� ��� �y�Դe�<����b��$�ԓ���%4����5�D�$���B{���-�� ����k6J���)��kZ�ۇk�tЪ�tU�S6���<m}��^�f+�,�+�u7r�@�;��o�&h������3��]b�/h�8�s7)t��_��E���h�������Df�/>�f�'����m�Q���?*@�$Y���<��$��[�X��A��DT��'	�.��c�),-~fMką4����Ħ)�oOi�p�=��ju�Y�ܪBu�qG�L�\����_�e�\}bm��yzE���s c�R�-	!N8��I�:�ڹ���]i���/=G��}EfOt-��[lX�	o��(�c@a�5`���������|zѩ�;^���&ѭ�kٱ|�Jiz�,�=~�!4�%17��~����2+5�B�����0Qהw0�-R��&���p)���5��WO�/4]��W�u��{/���!e`�/�Vށ�@�3D�n�6���͇��������է itE���\B�Wr���罯~�+����|����i�������V" ���`؛��KHt�\4Ԯ��I<>�83���)��g
��y-�dݾ�����2]�@ܘ�Y�������Ax(��" 7L�/F���_	F�U�@�OO���K�L��c�Qc�A���5�&-
�Nc Qu�"���8�V�{[:eF�9�v�\k�5yơ��F��N��^��d�/X/kU�u�k���Zȇq�a��&A�}�'p��� :}Q����H�`q�0��ȳ=�|T�tp1��!Dr�U�`�~dG6��l���}��g�$�"��%��	E'��d �8o_������6�2�r4���tlz�ٻ���<;eq;�TN�O����B�2C:-�d��I��\n�]�������V]�� �ǅ��4���m�r�x��"�7�@�g���V�P�+j%�	R���J�r;p��?�U��5h볅������x�D5�^�?}�i �c�?PD)���r�@��q��l�߶N�C�_��7N�E���Y���qc�s���/Q'p�(��
���X?X�_(G*��&w#ʮc!î��3�Tׄ\�e�Pa\�E��[TC/7F�a�li{ox ��<��6�J�Rz[73똗�ME�7��:C�~�
ư����CK��̈�E��Ճ�e:��ȁ������� �^������M�27��#za��SZ�9����7Y
��1� ����ۛe(߉]1�o�)^%��kj�Sm�P-�"�*V�j򮯝�#���km˖�؉�c��*+E���DT[e��PO�O�F��W�ʦHP�E�}!p��������'������C
*��JR�e��=�4�%���3X�M�M܆U���6/x+�����䖊�@�=�-�	ł滯���U��f ZL��8�+&�ˁ�d��������Q�70,V�U��X�½�4�3�)�a�(����p�]��
5��/��|%Y�]�W����]6~t{2��-��S(��G�ͧ�.��C��G���3┰r$o�#s�R��^��7�@CJ�S��K�Bs+�a»;-����p �j�KUAu���yU-N�sPv�'X"�	\�a�T�Sx4���w��pm��WE�}���2SU	1�O��I8�I���IN��wb�lG_��iӤ/�Th��A��E�M�4��YA�q�$�r���;'ΈW�q���aVM0��֋y怣�Yy\����-���t�h����p3���5�2���t�}V�����e�K^s�d�W�O��(��h\T#�j�F�
�U�eɘH�1����o�YS��V䮟�L���ޮ�H�v��;�KEW���<a�>����F��2�k��/n�s��Z"�:��*��[����
����s
�F+J�h{���[�DM�dL�=}��h\�4���ɍ=��ƌ����0N��'C����^��8q�����QS��(���񖿑|�y�5�-J>em�n�L1$V�����K*�%��!s>�WƤ��C ����g��,�(�v�+q)��J��R ;�ګ8]'7���|r(�m���Ҝ�7LЖ�w���]\�I���xHXPC<�����ip���������,�2jj��zδ��0*����n�F4ߛ�e�+��|��<]�l�=G����HW���x��m�E�sy�N�+I���X�\����C�`:xe��Q��2�ï*��[r�!)ifz.����J`7n<PI�}L͑J����e���f��5���0z>�)��L"��읙���њ�O�"�āu�&�#���d�n�m���L���jwo�ˉs;լ�����U��->o\Lf¸$�k��� !��L�bFK���C)u��k���>c��r�ѵV���P�-����"�̆ν���ty ����b$ɇT[�=��<ȫ��-+�Ӯ��-�#(DM*4Ǩ�&Bْ��Z�Bp@�>#P���"�������,����
�D#�0���{�8��c
�\���BF[?�z�Ѧ�;oMZCޒp#��+���&g�P��I13up��X�Ι�J���l��0V��Kw�~":�%# �P�eu=c$=��Ȟ�e	F��<��a��#z���i7-Xdq���i���]�s��c^�BNS"�-KB���~7G"���o+���:�QOϓy����yۤ30,H�Y��� +5�9Y��9����Ay�M{b��DCɸ��&�.sVИ�M�:����A��t������2�@��������uh�Y.�F��G�7-=7Ns�w�>ʊ�w� 2�=�j��[3RӴx´�{<���!��g���A���ӛ�/

Pg��5�#��7�fof��!�ǻm���i0���Ux�[Cz����[��4
S0��M� ��ft;�𱈮���n���y���'���*�wxޗ>���2�z��<ᄯZC�J��ꟶl���N��߫!+ƭ��&�q8͗	����أChR��#}Q=eW�Y�bһ�S�ҭ�<���蛜��)�4�,v� �W��m�5$�����]�E��m ��Gl4v@[�H�@��P��e����z�a�9����ƹ>ꌗ
s��`�Xs���i9�
�������]E���H�]n�&��G���8jX穚�q�x�����0Z�Lܒ�e���p��������c�H��iW`��!����"҂j2��p/5�� �in��t�ꫨh�=T�>�Sp���������p�*����Qs��E�D���o~�