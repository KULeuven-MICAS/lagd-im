// Copyright 2025 KU Leuven.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
// Author: Jiacong Sun <jiacong.sun@kuleuven.be>

`timescale 1ns / 1ps

`ifndef DBG
`define DBG 0
`endif

`ifndef VCD_FILE
`define VCD_FILE "tb_digital_macro.vcd"
`endif

`define True 1'b1
`define False 1'b0

`ifndef DataFromFile
`define DataFromFile `True
`endif

`ifndef EnComparison
`define EnComparison `True
`endif

`ifndef EnableFlipDetection
`define EnableFlipDetection `True
`endif

`ifndef FlipDisable
`define FlipDisable `True
`endif

`ifndef EnableAnalogLoop
`define EnableAnalogLoop `True
`endif

`ifndef MultiCmptModeEn
`define MultiCmptModeEn `False
`endif

module tb_digital_macro;
    import analog_format_pkg::*;
    import energy_calc_pkg::*;
    import config_pkg::*;
    import data_read_pkg::*;

    // testbench parameters
    localparam int CLKCYCLE = 2;
    localparam int NUM_TESTS = 1; // number of computation processes (only 1 is supported currently)

    // dut signals
    logic clk_i;
    logic rst_ni;
    logic en_aw_i, en_fm_i, en_em_i, en_ff_i, en_ef_i, en_analog_loop_i, en_perf_counter_i;
    logic en_i;
    logic config_valid_em_i;
    logic config_valid_fm_i;
    logic config_valid_aw_i;
    logic debug_dt_configure_enable_i;
    logic debug_spin_configure_enable_i;
    logic [ $clog2(NUM_SPIN)-1 : 0 ] config_counter_i;
    logic [ NUM_SPIN*SPIN_DEPTH-1 : 0 ] config_spin_initial_i;
    logic [ SPIN_DEPTH-1 : 0 ] config_spin_initial_skip_i;
    logic [ COUNTER_BITWIDTH-1 : 0] cfg_trans_num_i;
    logic [ COUNTER_BITWIDTH-1 : 0] cycle_per_wwl_high_i;
    logic [ COUNTER_BITWIDTH-1 : 0] cycle_per_wwl_low_i;
    logic [ COUNTER_BITWIDTH-1 : 0] cycle_per_spin_write_i;
    logic [ COUNTER_BITWIDTH-1 : 0] cycle_per_spin_compute_i;
    logic [ NUM_SPIN : 0 ] wwl_vdd_i;
    logic [ NUM_SPIN : 0 ] wwl_vread_i;
    logic [ NUM_SPIN : 0 ] wwl_vdd_o;
    logic [ NUM_SPIN : 0 ] wwl_vread_o;
    logic bypass_data_conversion_i;
    logic [ NUM_SPIN-1 : 0 ] spin_wwl_strobe_i;
    logic [ NUM_SPIN-1 : 0 ] spin_feedback_i;
    logic [ $clog2(SYNCHRONIZER_PIPEDEPTH)-1 : 0 ] synchronizer_pipe_num_i;
    logic [ $clog2(SYNCHRONIZER_PIPEDEPTH)-1 : 0 ] synchronizer_wbl_pipe_num_i;
    logic dt_cfg_enable_i, dt_cfg_idle_o;
    logic j_mem_ren_o;
    logic [ $clog2(NUM_SPIN / PARALLELISM)-1 : 0 ] j_raddr_o, dgt_weight_raddr_o;
    logic [ NUM_SPIN*BITJ*PARALLELISM-1 : 0 ] j_rdata_i, dgt_weight_i;
    logic h_ren_o;
    logic [ BITH*NUM_SPIN-1 : 0 ] h_rdata_i;
    logic flush_i;
    logic en_comparison_i;
    logic cmpt_en_i;
    logic cmpt_idle_o;
    logic host_readout_i;
    logic flip_ren_o;
    logic [ $clog2(FLIP_ICON_DEPTH)-1 : 0 ] flip_raddr_o, flip_raddr_ref;
    logic [ $clog2(FLIP_ICON_DEPTH)+1-1 : 0 ] icon_last_raddr_plus_one_i;
    logic [ NUM_SPIN-1 : 0 ] flip_rdata_i;
    logic flip_disable_i;
    logic [ BITH*NUM_SPIN-1 : 0 ] dgt_hbias_i;
    logic [ SCALING_BIT-1 : 0 ] dgt_hscaling_i;
    logic [ NUM_SPIN-1 : 0 ] j_one_hot_wwl_o;
    logic h_wwl_o;
    logic [NUM_SPIN*BITJ-1 : 0 ] wbl_o;
    logic [NUM_SPIN*BITJ-1 : 0 ] wblb_o;
    logic [NUM_SPIN*BITJ-1 : 0 ] wbl_floating_i, wbl_floating_o;
    logic [ NUM_SPIN-1 : 0 ] spin_wwl_o;
    logic [NUM_SPIN-1 : 0 ] spin_feedback_o;
    logic [ NUM_SPIN-1 : 0 ] spin_analog_i;
    logic signed [SPIN_DEPTH-1:0] [ENERGY_TOTAL_BIT-1:0] energy_fifo_o;
    logic [SPIN_DEPTH-1:0] [NUM_SPIN-1:0] spin_fifo_o;
    logic dgt_weight_ren_o;
    logic [ $clog2(NUM_SPIN / PARALLELISM)-1 : 0 ] dgt_addr_upper_bound_i;
    logic energy_fifo_update_o;
    logic spin_fifo_update_o;
    logic enable_flip_detection_i;
    logic debug_spin_compute_en_i;
    logic infinite_icon_loop_en_i;
    logic multi_cmpt_mode_en_i;
    logic [CC_COUNTER_BITWIDTH-1:0] cmpt_cycle_cnt_o;
    logic cmpt_cycle_cnt_maxed_o;
    logic cmpt_cycle_cnt_overflow_o;

    // debugging interface
    logic [COUNTER_BITWIDTH-1:0] debug_cycle_per_spin_read_i;
    logic [COUNTER_BITWIDTH-1:0] debug_spin_read_num_i;
    logic debug_j_write_en_i;
    logic debug_j_read_en_i;
    logic [NUM_SPIN-1:0] debug_j_one_hot_wwl_i;
    logic debug_h_wwl_i;
    logic [NUM_SPIN*BITDATA-1:0] debug_wbl_i;
    logic debug_spin_write_en_i;
    logic debug_spin_read_en_i;
    logic debug_spin_valid_o;
    logic [DEBUG_WADDR_WIDTH-1:0] debug_spin_waddr_o;
    logic [NUM_SPIN-1:0] debug_spin_o;
    logic debug_j_read_data_valid_o;
    logic [NUM_SPIN*BITDATA-1:0] debug_j_read_data_o;
    logic [NUM_SPIN*BITDATA-1:0] wbl_read_i, wblb_read_i;

    // testbench signals
    logic config_em_done;
    logic config_fm_done;
    logic config_aw_done;
    logic config_galena_done;
    logic config_dut_done;
    logic [ $clog2(NUM_SPIN / PARALLELISM)-1 : 0 ] j_raddr_ref, weight_raddr_ref;
    logic [NUM_SPIN*BITJ-1:0] wbl_copy;
    logic [NUM_SPIN-1:0][NUM_SPIN*BITJ-1:0] weights_in_txt, weights_analog;
    logic [NUM_SPIN/PARALLELISM-1:0][NUM_SPIN*BITJ*PARALLELISM-1:0] weights_in_mem;
    logic [NUM_SPIN*BITH-1:0] hbias_in_reg, hbias_analog;
    logic [SCALING_BIT-1:0] hscaling_in_reg;
    logic [SPIN_DEPTH-1:0] [NUM_SPIN-1:0] spin_initial_states;
    logic [NUM_SPIN*BITDATA-1:0] wbl_i;
    int signed constant;
    logic [IconLastAddrPlusOne-1:0] [NUM_SPIN-1:0] flip_icons_in_mem;
    logic signed [IconLastAddrPlusOne-1+1:0] [SPIN_DEPTH-1:0] [ENERGY_TOTAL_BIT-1:0] energy_fifo_ref;
    logic [IconLastAddrPlusOne-1+1:0] [SPIN_DEPTH-1:0] [NUM_SPIN-1:0] spin_fifo_ref;
    int unsigned total_cycles, transaction_cycles, total_time, transaction_time, start_time, end_time;
    int test_idx;
    logic cmpt_test_start, cmpt_test_end;
    logic final_fifo_check_end;
    integer dt_write_cycle_cnt_j;
    logic [IconLastAddrPlusOne-1:0] [NUM_SPIN-1:0] states_out_ref;
    model_t model_data;
    logic [CC_COUNTER_BITWIDTH-1:0] cmpt_max_num_i;
    logic multi_cmpt_mode_idle_o;
    logic [CC_COUNTER_BITWIDTH-1:0] cmpt_idx_o, cycle_per_iteration_o, cycle_per_cmpt_o;
    logic [2*CC_COUNTER_BITWIDTH-1:0] cycle_all_cmpt_o;
    logic [COUNTER_BITWIDTH-1:0] multi_cmpt_idx;

    assign en_aw_i = en_i;
    assign en_em_i = en_i;
    assign en_fm_i = en_i;
    assign en_ff_i = en_i;
    assign en_perf_counter_i = en_i;
    assign dgt_addr_upper_bound_i = NUM_SPIN / PARALLELISM - 1;
    assign debug_dt_configure_enable_i = 1'b0;
    assign debug_spin_configure_enable_i = 1'b0;
    assign wwl_vdd_i = {NUM_SPIN+1{1'b1}}; // all VDDs are enabled
    assign wwl_vread_i = {NUM_SPIN+1{1'b0}}; // all VREADs are disabled
    assign debug_cycle_per_spin_read_i = 'd0;
    assign debug_spin_read_num_i = 'd0;
    assign infinite_icon_loop_en_i = INFINITE_ICON_LOOP_EN;
    assign multi_cmpt_mode_en_i = `MultiCmptModeEn;
    assign cmpt_max_num_i = CmptMaxNum - 1; // max number of computations in multi-cmpt mode

    always_comb begin
        for (int i=0; i < NUM_SPIN; i=i+1) begin
            spin_analog_i[i] = wbl_i[i*BITDATA + SPIN_WBL_OFFSET];
        end
    end

    // module instantiation
    digital_macro #(
        .BITJ                            (BITJ                          ),
        .BITH                            (BITH                          ),
        .NUM_SPIN                        (NUM_SPIN                      ),
        .SCALING_BIT                     (SCALING_BIT                   ),
        .PARALLELISM                     (PARALLELISM                   ),
        .ENERGY_TOTAL_BIT                (ENERGY_TOTAL_BIT              ),
        .LITTLE_ENDIAN                   (LITTLE_ENDIAN                 ),
        .PIPESINTF                       (PIPESINTF                     ),
        .PIPESMID                        (PIPESMID                      ),
        .PIPESFLIPFILTER                 (PIPESFLIPFILTER               ),
        .SPIN_DEPTH                      (SPIN_DEPTH                    ),
        .FLIP_ICON_DEPTH                 (FLIP_ICON_DEPTH               ),
        .COUNTER_BITWIDTH                (COUNTER_BITWIDTH              ),
        .SYNCHRONIZER_PIPEDEPTH          (SYNCHRONIZER_PIPEDEPTH        ),
        .SPIN_WBL_OFFSET                 (SPIN_WBL_OFFSET               ),
        .H_IS_NEGATIVE                   (H_IS_NEGATIVE                 ),
        .ENABLE_FLIP_DETECTION           (ENABLE_FLIP_DETECTION         ),
        .CC_COUNTER_BITWIDTH             (CC_COUNTER_BITWIDTH           )
    ) dut (
        .clk_i                           (clk_i                         ),
        .rst_ni                          (rst_ni                        ),
        .en_aw_i                         (en_aw_i                       ),
        .en_em_i                         (en_em_i                       ),
        .en_ff_i                         (en_ff_i                       ),
        .en_fm_i                         (en_fm_i                       ),
        .en_ef_i                         (en_ef_i                       ),
        .en_analog_loop_i                (en_analog_loop_i              ),
        .en_perf_counter_i               (en_perf_counter_i             ),
        .config_valid_em_i               (config_valid_em_i             ),
        .config_valid_fm_i               (config_valid_fm_i             ),
        .config_valid_aw_i               (config_valid_aw_i             ),
        .debug_dt_configure_enable_i     (debug_dt_configure_enable_i   ),
        .debug_spin_configure_enable_i   (debug_spin_configure_enable_i ),
        .config_counter_i                (config_counter_i              ),
        .config_spin_initial_i           (config_spin_initial_i         ),
        .config_spin_initial_skip_i      (config_spin_initial_skip_i    ),
        .cfg_trans_num_i                 (cfg_trans_num_i               ),
        .cycle_per_wwl_high_i            (cycle_per_wwl_high_i          ),
        .cycle_per_wwl_low_i             (cycle_per_wwl_low_i           ),
        .cycle_per_spin_write_i          (cycle_per_spin_write_i        ),
        .cycle_per_spin_compute_i        (cycle_per_spin_compute_i      ),
        .wwl_vdd_i                       (wwl_vdd_i                     ),
        .wwl_vread_i                     (wwl_vread_i                   ),
        .bypass_data_conversion_i        (bypass_data_conversion_i      ),
        .spin_wwl_strobe_i               (spin_wwl_strobe_i             ),
        .spin_feedback_i                 (spin_feedback_i               ),
        .synchronizer_pipe_num_i         (synchronizer_pipe_num_i       ),
        .synchronizer_wbl_pipe_num_i     (synchronizer_wbl_pipe_num_i   ),
        .debug_cycle_per_spin_read_i     (debug_cycle_per_spin_read_i   ),
        .debug_spin_read_num_i           (debug_spin_read_num_i         ),
        .dt_cfg_enable_i                 (dt_cfg_enable_i               ),
        .j_mem_ren_o                     (j_mem_ren_o                   ),
        .j_raddr_o                       (j_raddr_o                     ),
        .j_rdata_i                       (j_rdata_i                     ),
        .h_ren_o                         (h_ren_o                       ),
        .h_rdata_i                       (h_rdata_i                     ),
        .dt_cfg_idle_o                   (dt_cfg_idle_o                 ),
        .flush_i                         (flush_i                       ),
        .en_comparison_i                 (en_comparison_i               ),
        .cmpt_en_i                       (cmpt_en_i                     ),
        .cmpt_idle_o                     (cmpt_idle_o                   ),
        .host_readout_i                  (host_readout_i                ),
        .flip_ren_o                      (flip_ren_o                    ),
        .flip_raddr_o                    (flip_raddr_o                  ),
        .icon_last_raddr_plus_one_i      (icon_last_raddr_plus_one_i    ),
        .flip_rdata_i                    (flip_rdata_i                  ),
        .flip_disable_i                  (flip_disable_i                ),
        .dgt_weight_ren_o                (dgt_weight_ren_o              ),
        .dgt_weight_raddr_o              (dgt_weight_raddr_o            ),
        .dgt_addr_upper_bound_i          (dgt_addr_upper_bound_i        ),
        .dgt_weight_i                    (dgt_weight_i                  ),
        .dgt_hbias_i                     (dgt_hbias_i                   ),
        .dgt_hscaling_i                  (dgt_hscaling_i                ),
        .j_one_hot_wwl_o                 (j_one_hot_wwl_o               ),
        .h_wwl_o                         (h_wwl_o                       ),
        .wbl_o                           (wbl_o                         ),
        .wblb_o                          (wblb_o                        ),
        .wbl_read_i                      (wbl_read_i                    ),
        .wblb_read_i                     (wblb_read_i                   ),
        .wbl_floating_o                  (wbl_floating_o                ),
        .wwl_vread_o                     (wwl_vread_o                   ),
        .wwl_vdd_o                       (wwl_vdd_o                     ),
        .spin_wwl_o                      (spin_wwl_o                    ),
        .spin_feedback_o                 (spin_feedback_o               ),
        .spin_analog_i                   (spin_analog_i                 ),
        .energy_fifo_update_o            (energy_fifo_update_o          ),
        .spin_fifo_update_o              (spin_fifo_update_o            ),
        .energy_fifo_o                   (energy_fifo_o                 ),
        .spin_fifo_o                     (spin_fifo_o                   ),
        .enable_flip_detection_i         (enable_flip_detection_i       ),
        // debugging interface
        .debug_j_write_en_i              (debug_j_write_en_i            ),
        .debug_j_read_en_i               (debug_j_read_en_i             ),
        .debug_j_one_hot_wwl_i           (debug_j_one_hot_wwl_i         ),
        .debug_h_wwl_i                   (debug_h_wwl_i                 ),
        .debug_wbl_i                     (debug_wbl_i                   ),
        .debug_j_read_data_o             (debug_j_read_data_o           ),
        .debug_j_read_data_valid_o       (debug_j_read_data_valid_o     ),
        .debug_spin_write_en_i           (debug_spin_write_en_i         ),
        .wbl_floating_i                  (wbl_floating_i                ),
        .debug_spin_compute_en_i         (debug_spin_compute_en_i       ),
        .debug_spin_read_en_i            (debug_spin_read_en_i          ),
        .debug_spin_valid_o              (debug_spin_valid_o            ),
        .debug_spin_waddr_o              (debug_spin_waddr_o            ),
        .debug_spin_o                    (debug_spin_o                  ),
        .debug_analog_dt_w_idle_o        (                              ),
        .debug_analog_dt_r_idle_o        (                              ),
        .debug_spin_w_idle_o             (                              ),
        .debug_spin_cmpt_idle_o          (                              ),
        .debug_spin_r_idle_o             (                              ),
        .debug_fm_upstream_handshake_o   (                              ),
        .debug_fm_energy_input_o         (                              ),
        .debug_fm_downstream_handshake_o (                              ),
        .debug_fm_spin_out_o             (                              ),
        .debug_aw_downstream_handshake_o (                              ),
        .debug_aw_spin_out_o             (                              ),
        .debug_em_upstream_handshake_o   (                              ),
        .debug_em_spin_in_o              (                              ),
        // measurement purposes
        .infinite_icon_loop_en_i         (infinite_icon_loop_en_i       ),
        .multi_cmpt_mode_en_i            (multi_cmpt_mode_en_i          ),
        .cmpt_max_num_i                  (cmpt_max_num_i                ),
        .multi_cmpt_mode_idle_o          (multi_cmpt_mode_idle_o        ),
        .cmpt_idx_o                      (cmpt_idx_o                    ),
        .cycle_per_iteration_o           (cycle_per_iteration_o         ),
        .cycle_per_cmpt_o                (cycle_per_cmpt_o              ),
        .cycle_all_cmpt_o                (cycle_all_cmpt_o              )
    );

    // Clock generation
    initial begin
        clk_i = 0;
        forever #(CLKCYCLE/2) clk_i = ~clk_i;
    end

    // Reset and en_i generation
    initial begin
        rst_ni = 0;
        en_i = 0;
        en_analog_loop_i = 0;
        #(5 * CLKCYCLE);
        rst_ni = 1;
        #(5 * CLKCYCLE);
        en_i = 1;
        en_analog_loop_i = `EnableAnalogLoop;
    end

    // Run tests
    initial begin
        if (`DBG) begin
            $display("Debug mode enabled. Running with detailed output.");
            $timeformat(-9, 1, " ns", 9);
            $dumpfile(`VCD_FILE);
            $dumpvars(1, tb_digital_macro); // Dump all variables in testbench module
            #(1000 * CLKCYCLE); // To avoid generating huge VCD files
            $display("[Time: %t] Testbench timeout reached. Ending simulation.", $time);
            $finish;
        end
        else begin
            $timeformat(-9, 1, " ns", 9);
            if (`MultiCmptModeEn) begin
                #(500_000 * CmptMaxNum * CLKCYCLE);
            end else begin
                #(500_000 * CLKCYCLE);
            end
            $display("[Time: %t] Testbench timeout reached. Ending simulation.", $time);
            $finish;
        end
    end

    initial begin
        en_ef_i = 0;
        wait (cmpt_en_i == 1);
        en_ef_i = 1;
        $display("[Time: %t] Energy monitor fifo starts to be enabled.", $time);
    end

    // ========================================================================
    // Functions
    // ========================================================================
    // Generate random model
    // note: the most negative code (-8), though supported by the digital logic, is not supported by the analog part and its related data convertor
    // therefore, we should avoid generating this code here
    function automatic model_t generate_random_model();
        model_t model;
        for (int i = 0; i < NUM_SPIN; i = i + 1) begin
            for (int j = 0; j < NUM_SPIN; j = j + 1) begin
                if (LITTLE_ENDIAN) begin
                    if (j == i) begin
                        model.weights[i][j*BITJ +: BITJ] = 'd0;
                    end else begin
                        do begin
                            model.weights[i][j*BITJ +: BITJ] = $urandom_range(0, (1<<BITJ)-1);
                        end while (model.weights[i][j*BITJ +: BITJ] == {1'b1, {BITJ-1{1'b0}}}); // avoid generating the invalid code
                    end
                end else begin
                    if (j == NUM_SPIN - 1 - i) begin
                        model.weights[i][j*BITJ +: BITJ] = 'd0;
                    end else begin
                        do begin
                            model.weights[i][j*BITJ +: BITJ] = $urandom_range(0, (1<<BITJ)-1);
                        end while (model.weights[i][j*BITJ +: BITJ] == {1'b1, {BITJ-1{1'b0}}}); // avoid generating the invalid code
                    end
                end
            end
        end
        // ensure matrix J is symmetric
        for (int i = 0; i < NUM_SPIN; i = i + 1) begin
            for (int j = i+1; j < NUM_SPIN; j = j + 1) begin
                if (LITTLE_ENDIAN) begin
                    model.weights[j][i*BITJ +: BITJ] = model.weights[i][j*BITJ +: BITJ];
                end else begin
                    model.weights[j][(NUM_SPIN-1 - i)*BITJ +: BITJ] = model.weights[i][(NUM_SPIN-1 - j)*BITJ +: BITJ];
                end
            end
        end
        // generate random h
        for (int i = 0; i < NUM_SPIN; i = i + 1) begin
            do begin
                model.hbias[i*BITH +: BITH] = $urandom_range(0, (1<<BITH)-1);
            end while (model.hbias[i*BITH +: BITH] == {1'b1, {BITH-1{1'b0}}}); // avoid generating the invalid code
        end
        // generate random scaling factor
        model.scaling_factor = $urandom_range(0, 2**SCALING_BIT-1);
        // constant
        model.constant = 0;
        return model;
    endfunction

    // ========================================================================
    // Sub-tasks
    // ========================================================================
    // Generate weight model
    task automatic gen_model();
        if (`DataFromFile == `False) begin: randomly_generate_model
            model_data = generate_random_model();
        end else begin: load_model_from_file
            model_data = load_model();
        end
        weights_in_txt = model_data.weights;
        hbias_in_reg = model_data.hbias;
        hscaling_in_reg = model_data.scaling_factor;
        constant = model_data.constant;

        // map to memory format
        for (int i = 0; i < NUM_SPIN/PARALLELISM; i = i + 1) begin
            for (int j = 0; j < PARALLELISM; j = j + 1) begin
                weights_in_mem[i][j*NUM_SPIN*BITJ +: NUM_SPIN*BITJ] = weights_in_txt[i*PARALLELISM + j];
            end
        end
    endtask

    // Generate flipping icons
    task automatic gen_flip_icons();
        if (`DataFromFile == `True) begin: load_flip_icons_from_file
            flip_icons_in_mem = load_flip_icons();
        end else begin: randomly_generate_flip_icons
            for (int i = 0; i < IconLastAddrPlusOne; i = i + 1) begin
                for (int j = 0; j < NUM_SPIN; j = j + 1) begin
                    flip_icons_in_mem[i][j] = $urandom_range(0, 1);
                end
            end
        end
    endtask

    // Generate initial spin states
    task automatic gen_initial_states();
        if (`DataFromFile == `True) begin: load_initial_states_from_file
            spin_initial_states = load_initial_states();
        end else begin: randomly_generate_initial_states
            for (int i = 0; i < SPIN_DEPTH; i = i + 1) begin
                for (int j = 0; j < NUM_SPIN; j = j + 1) begin
                    spin_initial_states[i][j] = $urandom_range(0, 1);
                end
            end
        end
    endtask

    // Generate reference model for spin fifo
    task automatic gen_ref_energy_spin_fifo();
        logic signed [ENERGY_TOTAL_BIT-1:0] energy_temp = 0;
        integer spin_fifo_pointer = 0;
        logic [NUM_SPIN-1:0] current_spin_state;

        if (`DataFromFile == `True && `EnableAnalogLoop == `True) begin
            states_out_ref = load_state_out_ref();
        end else begin
            states_out_ref = 'd0; // not used
        end

        for (int i = 0; i < SPIN_DEPTH; i = i + 1) begin
            spin_fifo_ref[0][i] = spin_initial_states[i];
            energy_fifo_ref[0][i] = {1'b0, {(ENERGY_TOTAL_BIT-1){1'b1}}};
        end

        for (int icon_idx = 1; icon_idx <= IconLastAddrPlusOne; icon_idx = icon_idx + 1) begin
            // get current spin state
            if (`DataFromFile == `True && `EnableAnalogLoop == `True) begin
                current_spin_state = states_out_ref[icon_idx-1];
            end else begin
                current_spin_state = `FlipDisable ? spin_fifo_ref[icon_idx-1][spin_fifo_pointer] :
                    spin_fifo_ref[icon_idx-1][spin_fifo_pointer] ^ flip_icons_in_mem[icon_idx-1];
            end
            // calc energy
            energy_temp = calculate_h_energy(
                current_spin_state,
                weights_in_txt,
                hbias_in_reg,
                hscaling_in_reg
            );
            // update fifo
            for (int j = 0; j < SPIN_DEPTH; j = j + 1) begin
                if (j != spin_fifo_pointer) begin
                    spin_fifo_ref[icon_idx][j] = spin_fifo_ref[icon_idx-1][j];
                    energy_fifo_ref[icon_idx][j] = energy_fifo_ref[icon_idx-1][j];
                end
            end
            if (`EnComparison == `False) begin: always_update_fifo
                energy_fifo_ref[icon_idx][spin_fifo_pointer] = energy_temp;
                spin_fifo_ref[icon_idx][spin_fifo_pointer] = current_spin_state;
            end else begin: conditional_update_fifo
                if (energy_temp < $signed(energy_fifo_ref[icon_idx-1][spin_fifo_pointer])) begin
                    energy_fifo_ref[icon_idx][spin_fifo_pointer] = energy_temp;
                    spin_fifo_ref[icon_idx][spin_fifo_pointer] = current_spin_state;
                end else begin
                    energy_fifo_ref[icon_idx][spin_fifo_pointer] = energy_fifo_ref[icon_idx-1][spin_fifo_pointer];
                    spin_fifo_ref[icon_idx][spin_fifo_pointer] = spin_fifo_ref[icon_idx-1][spin_fifo_pointer];
                end
            end
            // update pointer
            spin_fifo_pointer = (spin_fifo_pointer + 1) % SPIN_DEPTH;
        end
        if (`DataFromFile == `True) begin
            $display("[Time: %t] Reference energy and spin fifo loaded from file.", $time);
            // output energies and states to files
            output_energies_to_file(energy_fifo_ref, model_data.constant);
            output_spins_to_file(spin_fifo_ref);
            $display("[Time: %t] Reference energy and spin fifo output to files.", $time);
        end else begin
            $display("[Time: %t] Reference energy and spin fifo generated.", $time);
        end
    endtask

    // Sub-task for AW config interface
    task automatic aw_config_interface();
        wait (rst_ni == 0);
        config_aw_done = 0;
        config_valid_aw_i = 0;
        cfg_trans_num_i = 'd0;
        cycle_per_wwl_high_i = 'd0;
        cycle_per_spin_write_i = 'd0;
        cycle_per_spin_compute_i = 'd0;
        synchronizer_pipe_num_i = 'd0;
        spin_wwl_strobe_i = 'd0;
        spin_feedback_i = 'd0;
        bypass_data_conversion_i = BypassDataConversion;
        // Apply configuration
        wait (rst_ni == 1 && en_i == 1);
        @(posedge clk_i);
        // $display("[Time: %t] AW configuration starts.", $time);
        config_valid_aw_i = 1;
        cfg_trans_num_i = NUM_SPIN/PARALLELISM-1+1;
        cycle_per_wwl_high_i = CyclePerWwlHigh - 1;
        cycle_per_wwl_low_i = CyclePerWwlLow - 1;
        cycle_per_spin_write_i = CyclePerSpinWrite - 1;
        cycle_per_spin_compute_i = CyclePerSpinCompute - 1;
        synchronizer_pipe_num_i = SynchronizerPipeNum;
        synchronizer_wbl_pipe_num_i = SynchronizerPipeNum;
        spin_wwl_strobe_i = SpinWwlStrobe;
        spin_feedback_i = SpinFeedback;
        @(posedge clk_i);
        config_valid_aw_i = 0;
        config_aw_done = 1;
        $display("[Time: %t] AW configuration finished.", $time);
    endtask

    // Sub-task for EM config interface
    task automatic em_config_interface();
        wait (rst_ni == 0);
        config_em_done = 0;
        config_valid_em_i = 0;
        config_counter_i = 'd0;
        wait (rst_ni == 1 && en_i == 1 && config_aw_done == 1);
        @(posedge clk_i);
        // $display("[Time: %t] EM configuration starts.", $time);
        config_valid_em_i = 1;
        config_counter_i = EmCfgCounter;
        @(posedge clk_i);
        config_valid_em_i = 0;
        config_em_done = 1;
        $display("[Time: %t] EM configuration finished.", $time);
    endtask

    // Sub-task for FM config interface
    task automatic fm_config_interface();
        wait (rst_ni == 0);
        config_fm_done = 0;
        config_valid_fm_i = 0;
        config_spin_initial_i = 'd0;
        config_spin_initial_skip_i = 'd0;
        flush_i = Flush;
        en_comparison_i = `EnComparison;
        icon_last_raddr_plus_one_i = IconLastAddrPlusOne;
        flip_disable_i = `FlipDisable;
        enable_flip_detection_i = `EnableFlipDetection;
        wait (rst_ni == 1 && en_i == 1 && config_em_done == 1);
        @(posedge clk_i);
        // $display("[Time: %t] FM configuration starts.", $time);
        config_spin_initial_i = spin_initial_states;
        config_spin_initial_skip_i = 'd0;
        config_valid_fm_i = 1'b1;
        @(posedge clk_i);
        config_valid_fm_i = 0;
        config_fm_done = 1;
        $display("[Time: %t] FM configuration finished.", $time);
    endtask

    // Sub-task for galena config
    task automatic galena_config_interface();
        wait (rst_ni == 0);
        config_galena_done = 0;
        dt_cfg_enable_i = 0;
        wait (rst_ni == 1 && en_i == 1 && config_aw_done == 1 && config_em_done == 1 && config_fm_done == 1);
        @(posedge clk_i);
        $display("[Time: %t] Galena configuration starts.", $time);
        dt_cfg_enable_i = 1;
        @(posedge clk_i);
        dt_cfg_enable_i = 0;
        @(posedge clk_i);
        wait (dt_cfg_idle_o == 1);
        config_galena_done = 1;
        $display("[Time: %t] Galena configuration finished.", $time);
    endtask

    // Sub-task for monitoring config done
    task automatic monitor_config_done();
        wait (rst_ni == 0);
        config_dut_done = 0;
        wait (config_aw_done == 1 && config_em_done == 1 && config_fm_done == 1 && config_galena_done == 1);
        @(posedge clk_i);
        config_dut_done = 1;
        $display("[Time: %t] DUT configuration is done.", $time);
    endtask

    // ========================================================================
    // Tasks
    // ========================================================================
    // Pre-compute configuration
    task automatic pre_compute_config();
        fork
            gen_flip_icons(); // generate flipping icons
            gen_initial_states(); // generate initial spin states
            gen_model(); // generate weight model
            gen_ref_energy_spin_fifo(); // generate reference energy and spin fifo
            aw_config_interface(); // configure aw module
            em_config_interface(); // configure em module
            fm_config_interface(); // configure fm module
            galena_config_interface(); // configure galena module
            monitor_config_done(); // monitor if dut config is done
        join_none
    endtask

    // Interface: analog_wrap <-> galena spin wwl
    task automatic galena_spin_wwl_interface();
        integer galena_spin_write_cycle_cnt = 0;
        wait (rst_ni == 1 && en_i == 1 && config_galena_done == 1);
        forever begin
            @(posedge clk_i);
            if ($countbits(spin_wwl_o, '1) == NUM_SPIN) begin: timer_start
                if (galena_spin_write_cycle_cnt == -1) begin: spin_write_finished
                    galena_spin_write_cycle_cnt = galena_spin_write_cycle_cnt;
                end else begin
                    if (galena_spin_write_cycle_cnt == (CyclePerSpinWrite-1)) begin: spin_write_finishing
                        wbl_copy = wbl_o;
                        galena_spin_write_cycle_cnt = -1;
                    end else begin: spin_write_ongoing
                        galena_spin_write_cycle_cnt = galena_spin_write_cycle_cnt + 1;
                    end
                end
            end else begin: spin_wwl_idle
                galena_spin_write_cycle_cnt = 0;
            end
        end
    endtask

    // Interface: analog_wrap <-> galena output
    task automatic galena_spin_output_interface();
        integer galena_spin_cmpt_cycle_cnt = 0;
        integer state_out_ref_idx = 0;

        wbl_i = 'd0;
        wait (rst_ni == 1 && en_i == 1 && config_galena_done == 1);
        forever begin
            @(posedge clk_i);
            wbl_i = 'z;
            if ($countbits(spin_wwl_o, '1) == NUM_SPIN) begin: timer_start
                while (galena_spin_cmpt_cycle_cnt < (CyclePerSpinWrite+CyclePerSpinCompute-2)) begin
                    galena_spin_cmpt_cycle_cnt = galena_spin_cmpt_cycle_cnt + 1;
                    if (galena_spin_cmpt_cycle_cnt >= CyclePerSpinWrite) begin
                        // during compute cycles, generate random wbl_i
                        for (int i = 0; i < NUM_SPIN * BITDATA; i = i + 1) begin
                            wbl_i[i] = $urandom_range(0, 1);
                        end
                    end
                    @(posedge clk_i);
                end
                // after compute cycles, output wbl_i
                if (`DataFromFile == `True) begin
                    for (int k = 0; k < NUM_SPIN; k = k + 1) begin
                        wbl_i[k*BITDATA] = {{(BITJ-1){1'b0}}, states_out_ref[state_out_ref_idx][k]} << SPIN_WBL_OFFSET;
                    end
                    state_out_ref_idx = (state_out_ref_idx + 1) % (IconLastAddrPlusOne);
                end else begin
                    wbl_i = wbl_copy;
                end
                galena_spin_cmpt_cycle_cnt = 0;
            end
        end
    endtask

    // Interface: J mem <-> analog wrap and energy monitor
    task automatic j_mem_interface();
        j_rdata_i = 'd0;
        dgt_weight_i = 'd0;
        j_raddr_ref = 'd0;
        weight_raddr_ref = 'd0;
        wait (rst_ni == 1 && en_i == 1);
        @(posedge clk_i);
        forever begin
            @(posedge clk_i);
            // Interface to analog wrap: standard 1-cycle-delay memory interface
            if (j_mem_ren_o == 1) begin
                if (j_raddr_o != j_raddr_ref) begin
                    $fatal(1, "[Time: %t] Error: J memory read address mismatch. Expected: %0d, Got: %0d",
                        $time, j_raddr_ref, j_raddr_o);
                end
                j_rdata_i = weights_in_mem[j_raddr_o];
                j_raddr_ref = j_raddr_ref + 1;
            end
            // Interface to energy monitor: standard 1-cycle-delay memory interface
            if (dgt_weight_ren_o == 1) begin
                if (ENABLE_FLIP_DETECTION == `False) begin
                    if (dgt_weight_raddr_o != weight_raddr_ref) begin
                        $fatal(1, "[Time: %t] Error: Weight memory read address mismatch. Expected: 'h%0h, Got: 'h%0h",
                            $time, weight_raddr_ref, dgt_weight_raddr_o);
                    end
                    dgt_weight_i = weights_in_mem[dgt_weight_raddr_o];
                    weight_raddr_ref = weight_raddr_ref + 1;
                end else begin
                    dgt_weight_i = weights_in_mem[dgt_weight_raddr_o];
                    weight_raddr_ref = dgt_weight_raddr_o + 1;
                end
            end
        end
    endtask

    // H and scaling factor reg interface
    task automatic h_sfc_reg_interface();
        h_rdata_i = hbias_in_reg; // for analog onloading
        dgt_hbias_i = hbias_in_reg; // for digital energy monitor
        dgt_hscaling_i = hscaling_in_reg;
    endtask

    // Flip icon memory interface
    task automatic flip_mem_interface();
        flip_rdata_i = 'd0;
        flip_raddr_ref = 'd0;
        wait (rst_ni == 1 && en_i == 1 && config_dut_done == 1);
        forever begin
            @(posedge clk_i);
            if (flip_ren_o == 1) begin
                if (flip_raddr_o != flip_raddr_ref) begin
                    $fatal(1, "[Time: %t] Error: Flip icon memory read address mismatch. Expected: %0d, Got: %0d",
                        $time, flip_raddr_ref, flip_raddr_o);
                end
                flip_rdata_i = flip_icons_in_mem[flip_raddr_o];
                flip_raddr_ref = flip_raddr_ref + 1;
            end
        end
    endtask

    // Host interface
    task automatic host_interface();
        host_readout_i = 0;
        test_idx = 0;
        cmpt_en_i = 0;
        cmpt_test_start = 0;
        cmpt_test_end = 0;
        wait (rst_ni == 1 && en_i == 1 && config_dut_done == 1);
        @(posedge clk_i);
        cmpt_test_start = 1;
        cmpt_en_i = 1;
        @(posedge clk_i);
        repeat (2) @(posedge clk_i);
        wait (final_fifo_check_end == 1);
        @(posedge clk_i);
        cmpt_test_end = 1;
    endtask

    // ========================================================================
    // Debug
    // ========================================================================
    task automatic debug_model_wr();
        debug_j_write_en_i = 1'b0;
        debug_j_read_en_i = 1'b0;
        debug_j_one_hot_wwl_i = 'd0;
        debug_h_wwl_i = 1'b0;
        debug_wbl_i = 'd0;
        wbl_floating_i = {(NUM_SPIN*BITDATA){1'b0}};
    endtask

    task automatic debug_model_spin_wr();
        debug_spin_write_en_i = 1'b0;
        debug_spin_read_en_i = 1'b0;
        debug_spin_compute_en_i = 1'b0;
    endtask

    // ========================================================================
    // Checks
    // ========================================================================
    // Task for analog galena interface: config data check: j
    task automatic analog_interface_config_check_j();
        integer config_test_correct_cnt_j = 0;
        integer galena_addr_idx = 0;
        dt_write_cycle_cnt_j = 0;
        while (config_test_correct_cnt_j < 1) begin
            wait (dt_cfg_enable_i == 1);
            @(posedge clk_i);
            // check if j and h are loaded correctly
            while (galena_addr_idx < NUM_SPIN) begin
                wait (j_one_hot_wwl_o != 0);
                while (dt_write_cycle_cnt_j < CyclePerWwlHigh) begin
                    @(negedge clk_i);
                    // monitor if j_one_hot_wwl_o remains valid for the dedefined cycles
                    if (j_one_hot_wwl_o == 0 && dt_write_cycle_cnt_j != 0) begin
                        $fatal(1, "[Time: %t] Warning: j_one_hot_wwl_o switches to zero during dt write cycle %0d for galena_addr_idx %0d",
                            $time, dt_write_cycle_cnt_j, galena_addr_idx);
                    end
                    if (|j_one_hot_wwl_o) begin
                        // check if one-hot encoded and matches galena_addr_idx
                        if ($countbits(j_one_hot_wwl_o, '1) != 1)
                            $fatal(1, "[Time: %t] Error: j_one_hot_wwl_o is not one-hot encoded, j_one_hot_wwl_o: 'b%b", $time, j_one_hot_wwl_o);
                        if (j_one_hot_wwl_o[galena_addr_idx] != 1'b1) begin
                            $fatal(1, "[Time: %t] Error: j_one_hot_wwl_o does not match galena_addr_idx, j_one_hot_wwl_o: 'b%b, galena_addr_idx: 'd%0d",
                                $time, j_one_hot_wwl_o, galena_addr_idx);
                        end
                        dt_write_cycle_cnt_j = dt_write_cycle_cnt_j + 1;
                    end
                end
                for (int i=0; i<NUM_SPIN; i=i+1) begin
                    if (bypass_data_conversion_i) begin: exact_copy_of_analog_data
                        weights_analog[galena_addr_idx][i*BITDATA +: BITDATA]
                            = wbl_o[i*BITDATA +: BITDATA];
                    end else begin: convert_data_format_for_checker
                        weights_analog[galena_addr_idx][i*BITDATA +: BITDATA]
                            = analog_to_signed_int(wbl_o[i*BITDATA +: BITDATA]);
                    end
                end
                // compare data to reference
                if (weights_analog[galena_addr_idx] != weights_in_txt[galena_addr_idx]) begin
                    $fatal(1, "[Time: %t] Error: Weights mismatch at galena_addr_idx %0d. Expected: 'h%h, Got: 'h%h",
                        $time, galena_addr_idx, weights_in_txt[galena_addr_idx], weights_analog[galena_addr_idx]);
                end
                dt_write_cycle_cnt_j = 0;
                galena_addr_idx = galena_addr_idx + 1;
            end
            config_test_correct_cnt_j = config_test_correct_cnt_j + 1;
            galena_addr_idx = 0;
        end
        // after all config tests
        $display("----------------------------------------");
        $display("Config Scoreboard [Time %0d ns]: %0d/%0d correct, %0d/%0d errors",
            $time, config_test_correct_cnt_j, 1, 1 - config_test_correct_cnt_j, 1);
        $display("----------------------------------------");
    endtask

    // Task for analog galena interface: config data check: h
    task automatic analog_interface_config_check_h();
        integer dt_write_cycle_cnt_hbias = 0;
        integer config_test_correct_cnt_h = 0;
        while (config_test_correct_cnt_h < 1) begin
            wait (rst_ni == 1 && en_i == 1);
            dt_write_cycle_cnt_hbias = 0;
            wait (dt_cfg_enable_i == 1);
            while (dt_write_cycle_cnt_hbias <  CyclePerWwlHigh) begin
                @(negedge clk_i);
                // monitor if h_wwl_o remains valid for the dedefined cycles
                if (h_wwl_o == 0 && dt_write_cycle_cnt_hbias != 0) begin
                    $fatal(1, "[Time: %t] Warning: h_wwl_o switches to zero during dt write cycle %0d for hbias",
                        $time, dt_write_cycle_cnt_hbias);
                end
                if (h_wwl_o == 1) begin
                    dt_write_cycle_cnt_hbias = dt_write_cycle_cnt_hbias + 1;
                end
            end
            // after dt write cycles, check hbias
            for (int i=0; i<NUM_SPIN; i=i+1) begin
                if (bypass_data_conversion_i) begin
                    hbias_analog[i*BITDATA +: BITDATA]
                    = wbl_o[i*BITDATA +: BITDATA];
                end else begin
                    hbias_analog[i*BITDATA +: BITDATA]
                        = analog_to_signed_int(wbl_o[i*BITDATA +: BITDATA]);
                end
            end
            // compare data to reference
            if (hbias_analog != hbias_in_reg) begin
                $fatal(1, "[Time: %t] Error: Hbias mismatch. Expected: 'h%h, Got: 'h%h",
                    $time, hbias_in_reg, hbias_analog);
            end
            config_test_correct_cnt_h = config_test_correct_cnt_h + 1;
        end
    endtask

    // Task for spin_wwl_o check
    task automatic spin_wwl_check();
        integer spin_wwl_cycle_cnt;
        spin_wwl_cycle_cnt = 0;
        wait (rst_ni == 1 && en_i == 1 && config_galena_done == 1);
        @(negedge clk_i);
        forever begin
            @(negedge clk_i);
            if ($countbits(spin_wwl_o, '1) != 0) begin
                if ($countbits(spin_wwl_o, '1) != NUM_SPIN) begin
                    $fatal(1, "[Time: %t] Error: spin_wwl_o is not all-one when enabled, spin_wwl_o: 'b%b",
                        $time, spin_wwl_o);
                end
                while (spin_wwl_cycle_cnt < CyclePerSpinWrite) begin
                    if (spin_wwl_cycle_cnt > 0 && $countbits(spin_wwl_o, '1) != NUM_SPIN) begin
                        $fatal(1, "[Time: %t] Error: spin_wwl_o is not all-one during spin write cycle %0d, spin_wwl_o: 'b%b",
                            $time, spin_wwl_cycle_cnt, spin_wwl_o);
                    end
                    spin_wwl_cycle_cnt = spin_wwl_cycle_cnt + 1;
                    @(negedge clk_i);
                end
                spin_wwl_cycle_cnt = 0;
            end
        end
    endtask

    // Check energy fifo content
    task automatic energy_fifo_check();
        integer test_correct_cnt = 0;
        integer check_idx = 0;

        multi_cmpt_idx = 0;
        wait (cmpt_test_start == 1);
        do begin
            check_idx = 0;
            test_correct_cnt = 0;
            while (check_idx < IconLastAddrPlusOne) begin
                while (energy_fifo_update_o == 0) @(negedge clk_i);
                for (int depth_idx = 0; depth_idx < SPIN_DEPTH; depth_idx = depth_idx + 1) begin
                    // check energy fifo
                    if (energy_fifo_o[depth_idx] !== energy_fifo_ref[check_idx+1][depth_idx]) begin
                        $fatal(1, "[Time: %t] Error: Energy fifo mismatch at check_idx 'd%0d, depth_idx 'd%0d. Expected: 'h%h, Got: 'h%h, hbias: 'h%h, hscaling: 'h%h, spin: 'h%h, state_out_ref: 'h%h",
                            $time, check_idx, depth_idx, energy_fifo_ref[check_idx+1][depth_idx], energy_fifo_o[depth_idx], hbias_in_reg, hscaling_in_reg, spin_fifo_ref[check_idx+1][depth_idx], states_out_ref[check_idx]);
                    end else begin
                        // $display("[Time: %t] Energy fifo match at check_idx 'd%0d, depth_idx 'd%0d. Value: 'h%h",
                        //     $time, check_idx, depth_idx, energy_fifo_o[depth_idx]);
                    end
                end
                test_correct_cnt = test_correct_cnt + 1;
                check_idx = check_idx + 1;
                @(negedge clk_i);
            end
            multi_cmpt_idx = multi_cmpt_idx + 1;
        end while (`MultiCmptModeEn && multi_cmpt_idx < CmptMaxNum);
        // after all tests
        if (`MultiCmptModeEn) begin
            $display("----------------------------------------");
            $display("Energy FIFO Scoreboard [Time %0d ns]: %0d/%0d correct, %0d/%0d errors, multi_cmpt_idx: %0d/%0d",
                $time, test_correct_cnt, IconLastAddrPlusOne, IconLastAddrPlusOne - test_correct_cnt, IconLastAddrPlusOne, multi_cmpt_idx, CmptMaxNum);
            $display("----------------------------------------");
        end else begin
            $display("----------------------------------------");
            $display("Energy FIFO Scoreboard [Time %0d ns]: %0d/%0d correct, %0d/%0d errors",
                $time, test_correct_cnt, IconLastAddrPlusOne, IconLastAddrPlusOne - test_correct_cnt, IconLastAddrPlusOne);
            $display("----------------------------------------");
        end
    endtask

    // Check spin fifo content
    task automatic spin_fifo_check();
        integer test_correct_cnt = 0;
        integer check_idx = 0;
        integer multi_spin_check_idx = 0;

        wait (cmpt_test_start == 1);
        do begin
            check_idx = 0;
            test_correct_cnt = 0;
            wait (dut.cmpt_en_fm == 1'b1); // wait for compute start
            repeat (2) @(posedge clk_i);
            while (check_idx < IconLastAddrPlusOne) begin
                while (spin_fifo_update_o == 0) @(negedge clk_i);
                for (int depth_idx = 0; depth_idx < SPIN_DEPTH; depth_idx = depth_idx + 1) begin
                    // check spin fifo
                    if (spin_fifo_o[depth_idx] !== spin_fifo_ref[check_idx+1][depth_idx]) begin
                        $fatal(1, "[Time: %t] Error: Spin fifo mismatch at check_idx 'd%0d, depth_idx 'd%0d. Expected: 'h%h, Got: 'h%h",
                            $time, check_idx, depth_idx, spin_fifo_ref[check_idx+1][depth_idx], spin_fifo_o[depth_idx]);
                    end else begin
                        // $display("[Time: %t] Spin fifo match at check_idx 'd%0d, depth_idx 'd%0d. Value: 'b%b",
                        //     $time, check_idx, depth_idx, spin_fifo_o[depth_idx]);
                    end
                end
                test_correct_cnt = test_correct_cnt + 1;
                check_idx = check_idx + 1;
                @(negedge clk_i);
            end
            multi_spin_check_idx = multi_spin_check_idx + 1;
        end while (`MultiCmptModeEn && multi_spin_check_idx < CmptMaxNum);
        // after all tests
        if (`MultiCmptModeEn) begin
            $display("----------------------------------------");
            $display("Spin FIFO Scoreboard [Time %0d ns]: %0d/%0d correct, %0d/%0d errors, multi_spin_check_idx: %0d/%0d",
                $time, test_correct_cnt, IconLastAddrPlusOne, IconLastAddrPlusOne - test_correct_cnt, IconLastAddrPlusOne, multi_spin_check_idx, CmptMaxNum);
            $display("----------------------------------------");
        end else begin
            $display("----------------------------------------");
            $display("Spin FIFO Scoreboard [Time %0d ns]: %0d/%0d correct, %0d/%0d errors",
                $time, test_correct_cnt, IconLastAddrPlusOne, IconLastAddrPlusOne - test_correct_cnt, IconLastAddrPlusOne);
            $display("----------------------------------------");
        end
    endtask

    // Host readout check
    task automatic host_readout_check();
        integer check_fifo_idx = 0;
        integer multi_final_check_idx = 0;

        final_fifo_check_end = 0;

        do begin
            wait (cmpt_idle_o == 0); // wait for compute start
            wait (cmpt_idle_o == 1); // wait for compute end
            @(negedge clk_i);
            while(check_fifo_idx < SPIN_DEPTH) begin
                if (`FlipDisable == `False) begin
                    if (spin_fifo_o[check_fifo_idx] !== spin_fifo_ref[IconLastAddrPlusOne][check_fifo_idx]) begin
                        $fatal(1, "[Time: %t] Error: Final spin fifo mismatch at test_idx 'd%0d, check_fifo_idx 'd%0d. Expected: 'h%0h, Got: 'h%0h",
                            $time, test_idx, check_fifo_idx, spin_fifo_ref[IconLastAddrPlusOne][check_fifo_idx], spin_fifo_o[check_fifo_idx]);
                    end
                end else begin
                    if (spin_fifo_o[check_fifo_idx] !== spin_fifo_ref[2][check_fifo_idx]) begin
                        $fatal(1, "[Time: %t] Error: Final spin fifo mismatch at test_idx 'd%0d, check_fifo_idx 'd%0d. Expected: 'h%0h, Got: 'h%0h",
                            $time, test_idx, check_fifo_idx, spin_fifo_ref[2][check_fifo_idx], spin_fifo_o[check_fifo_idx]);
                    end
                end
                // $display("[Time: %t] Final spin fifo check successfully at idx 'd%0d, value: 'b%0b",
                //     $time, check_fifo_idx, spin_fifo_o[check_fifo_idx]);
                if (`FlipDisable == `False) begin
                    if (energy_fifo_o[check_fifo_idx] !== energy_fifo_ref[IconLastAddrPlusOne][check_fifo_idx]) begin
                        $fatal(1, "[Time: %t] Error: Final energy fifo mismatch at test_idx 'd%0d, check_fifo_idx 'd%0d. Expected: 'h%h, Got: 'h%h",
                            $time, test_idx, check_fifo_idx, energy_fifo_ref[IconLastAddrPlusOne][check_fifo_idx], energy_fifo_o[check_fifo_idx]);
                    end
                end else begin
                    if (energy_fifo_o[check_fifo_idx] !== energy_fifo_ref[2][check_fifo_idx]) begin
                        $fatal(1, "[Time: %t] Error: Final energy fifo mismatch at test_idx 'd%0d, check_fifo_idx 'd%0d. Expected: 'h%h, Got: 'h%h",
                            $time, test_idx, check_fifo_idx, energy_fifo_ref[2][check_fifo_idx], energy_fifo_o[check_fifo_idx]);
                    end
                end
                // $display("[Time: %t] Final energy fifo check successfully at idx 'd%0d, value: 'h%h",
                //     $time, check_fifo_idx, energy_fifo_o[check_fifo_idx]);
                check_fifo_idx = check_fifo_idx + 1;
            end
            multi_final_check_idx = multi_final_check_idx + 1;
            check_fifo_idx = 0;
        end while (`MultiCmptModeEn && multi_final_check_idx < CmptMaxNum);
        final_fifo_check_end = 1;
    endtask

    // Multiple computation mode check
    task automatic multi_cmpt_idx_check();
        integer multi_cmpt_idx = 0;
        do begin
            wait (cmpt_idle_o == 0); // wait for compute start
            wait (cmpt_idle_o == 1); // wait for compute end
            if (`MultiCmptModeEn && cmpt_idx_o != multi_cmpt_idx) begin
                $fatal(1, "[Time: %t] Error: cmpt_idx_o mismatch in multiple computation mode. Expected: %0d, Got: %0d",
                    $time, multi_cmpt_idx, cmpt_idx_o);
            end
            multi_cmpt_idx = multi_cmpt_idx + 1;
        end while (`MultiCmptModeEn && multi_cmpt_idx < CmptMaxNum);
    endtask

    // Cmpt enable and timer
    task automatic cmpt_enable_and_timer();
        integer multi_cmpt_timer_idx = 0;
        wait (rst_ni == 0);
        total_cycles = 0;
        transaction_cycles = 0;
        total_time = 0;
        transaction_time = 0;
        start_time = 0;
        end_time = 0;
        wait (cmpt_test_start == 1);
        do begin
            wait (cmpt_idle_o == 0);
            start_time = $time;
            @(posedge clk_i);
            wait (cmpt_idle_o == 1);
            end_time = $time;
            // calculate compute cycles
            total_time = end_time - start_time;
            total_cycles = total_time / CLKCYCLE;
            transaction_cycles = total_cycles / IconLastAddrPlusOne;
            transaction_time = transaction_cycles * CLKCYCLE;
            $display("@@@@@@ Timer per Computation @@@@@@@@@@@@");
            $display("Timer [Time %0d ns]: start time: %0d ns, end time: %0d ns, duration: %0d ns, flips: %0d",
                $time, start_time, end_time, total_time, IconLastAddrPlusOne);
            $display("Timer [Time %0d ns]: Total cycles: %0d cc [%0d ns], Cycles/flip: %0d cc [%0d ns]",
                $time, total_cycles, total_time, transaction_cycles, transaction_time);
            $display("Timer [Time %0d ns]: MultiCmptModeEn: %d, multi_cmpt_timer_idx: %0d/%0d",
                $time, `MultiCmptModeEn, multi_cmpt_timer_idx, CmptMaxNum);
            $display("@@@@@@ Timer per Computation @@@@@@@@@@@@");
            multi_cmpt_timer_idx = multi_cmpt_timer_idx + 1;
        end while (`MultiCmptModeEn && multi_cmpt_timer_idx < CmptMaxNum);
        $finish;
    endtask

    // Task for timing record on each computation
    task automatic timing_record();
        logic [IconLastAddrPlusOne-1:0][31:0] cycle_cnt;
        integer idx = 0;
        integer time_a, time_b;

        wait (cmpt_en_i == 1);
        while (idx < IconLastAddrPlusOne) begin
            @(posedge clk_i);
            time_a = $time;
            wait (dut.fm_upstream_handshake == 1);
            @(posedge clk_i);
            time_b = $time;
            cycle_cnt[idx] = (time_b - time_a) / CLKCYCLE;
            // $display("[Time: %t] Timing record for icon idx %0d: %0d cycles", $time, idx, cycle_cnt[idx]);
            idx = idx + 1;
        end
        output_timing_record_to_file(cycle_cnt);

    endtask

    // ========================================================================
    // Event execution
    // ========================================================================
    initial begin
        fork
            pre_compute_config(); // configure aw, em, fm modules
            // interfaces
            galena_spin_wwl_interface();
            host_interface();
            galena_spin_output_interface();
            j_mem_interface();
            h_sfc_reg_interface();
            flip_mem_interface();
            // checks
            analog_interface_config_check_j();
            analog_interface_config_check_h();
            spin_wwl_check();
            energy_fifo_check();
            spin_fifo_check();
            host_readout_check();
            multi_cmpt_idx_check();
            // timer
            cmpt_enable_and_timer();
            timing_record();
            // debug
            debug_model_wr(); // inactive
            debug_model_spin_wr(); // inactive
        join_none
    end

endmodule
