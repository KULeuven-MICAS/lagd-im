// Copyright 2025 KU Leuven.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Author: Giuseppe Sarda <giuseppe.sarda@esat.kuleuven.be>

// User configuration for LAGD system

`ifndef LAGD_CONFIG_SVH
`define LAGD_CONFIG_SVH

    // Number of Ising cores in the system
    // Maximum is 14 (because of AXI ID width limitations)
    `ifndef NUM_ISING_CORES
        `define NUM_ISING_CORES 1
    `endif

    `ifndef L1_J_MEM_SIZE_B
        `define L1_J_MEM_SIZE_B 32*1024
    `endif

    `ifndef L1_H_MEM_SIZE_B
        `define L1_H_MEM_SIZE_B 128
    `endif

    `ifndef L1_FLIP_MEM_SIZE_B
        `define L1_FLIP_MEM_SIZE_B 32*1024
    `endif

    `ifndef L2_MEM_SIZE_B
        `define L2_MEM_SIZE_B 64*1024
    `endif

    `ifndef NUM_SPIN
        `define NUM_SPIN 256
    `endif

`endif // LAGD_CONFIG_SVH
