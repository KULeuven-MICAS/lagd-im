 GITCRYPT ��l9[}��W��ؠ�.44�"��"���A��|�M�J>�1^��Bn��ϥ(�3T�KU�c�vYx��k��X������S��=��=2l�B�f�vK�ʿB�n����fj�4��C��V3�)gT��.�1��C����Ax��C _[�	�r� r�2)8j!X���\u�6�n��E���Vh��?+0��
�����S2�#�:�r�g(Y�vϹ��BI �	�X���A�]��޾�x\h���M�3Hb�oK�z8�\��j��Xq���,t1��&>y
�b��.��d�KTҼL�8t�ߐ�>�1^/�l��115���"�^�I�@\� '����^����π�ji�"8/S��U�=�%�n�G{�#!ۈ�-ڷa�MoZ,� � <>`tv�C�1z���"o�1����Ѕ�6������E$�Ҩ�����`�^�+�>C��3ZD�aW�("VoV���u4���k�[�����M$��~�;a`2ލkk�u�)��K���^��X�g��?"��{{��7��	��J� .�!@|[�,�̱!��o��1)����/�d3{khA�_�Ϩ	N8O�\l����4S��q�^�V(��c)o=�t����QӨ��m�n���<�Uy���A?�3tN���I�`*vG�	O�&Y5@�:�kP��ʄ�I!g��=�C��XZ�F	��Zr�Ԉ�F �B,�OZ�5c�è�;j�e�1J 3������V-TX3�,�~7����t���i�%������XЋ�:�j�C7�����O�gBz�h+c5p~n�����)��t�E�AFcπ�YJQR��&���y��m��*��8�ۇ+��^"�'��{.ld����ي{�peϚ��y�Q=�B���x-C�BN�1L�t)���|��<K�SL $��@Ӏ�;�m��뒿��+\�|R�L�K�tD�P�Bly�?ZcLⰟ��bt�����ן-�窺��B� �p.��`D\�,�����n/86����٢؟��U������t�4����y���X���R~)�e�N���`�,ݝS�X&~����2��T��$�;�
�쥋$�E ���x�@���a�0���.�is�v��1b!v���:(g��(G��ΗV�8��hM�I�]�{�-%nM�UH�j_\rg��~#�۩�\x\3�a~-Z�� ̰��
�dU�y3<3pq �P��[�+S���?C�z�T��<������\ND�/��P�j����k`5����&1�; ��aJ�8�_��~N����՞|G�E�
��-�޼�p�^*ڄ�9���fҎ4�]�<��t��ֺ�?��uV�B��a�~IA����~�A)�3'uT/�ӻ��ۡv:>@ W�7�o�^��t�G	��Io��ǋ<�Fg��!�o��`:i��[*$���M�\[+<�ʨ+G4��"3on�	��T��iM�4�=r?��IvӞ�g�`~��!0�ܗA=�B/�t��L���/���s���j
���)X��|���҂�`����`����˛o=>��7�=��L�K�کp����^������-z���BEp�#��8N��\��(+o�J�H�ͅI�I1i�*3��������єva��ע�*^��M�|X�F8ͩMŊ��T�RA��Ծ���kd}��4׃`OR�'��s��z]���UY���򇖻_�I"�oL�\�/�_�Xu�{	8N�N�p(���0�a��Ā+�!{;�lmS�!ME�%df�Lߧ��mw^���j�`����),U[�)N����d�)�[��,SK������AN]������t�utZ����g^�H.	u��f/�����,�2!m������7-1��F3��2l���ڜ�.�]y����J�2(�8�'�{P�j�����W�<������(���	����RJH��{
	�(�F�-���O�aX����Ќ)�tI�d4�d�� ��ӕ�w����A�au�ؒ��gԏ�-\�҃g�X8�T80�d�/_6.m�d�$����g�J�~wB�̓�x>���DH�VKU���[�a���i��-緪g�B:Y5��s��C6�e��4��}q�!Z=`[��[��		hN��D��:�C�}�Ξ���A�%{3�s��x2:�����㐋� ���bq>�_[	��%9"���I�V��
��v_A���n�8�9"��P�N�ق��v� �&���a�bm�x'9���HsOk��nR�(��5SF��!��*Ɓ�@_��0�b)�����I^���lMRC���q��1i�R�nO�@�\rH�ۺ�h�E��<� �T�����j�Or	7�(@^��̀���DG�]\lg��;{�XQ�����U��A�����J8ݗ*>y���IFӏ�E���Dk�?�y�T���+H���1H���T,�m���M�)�72��ϾTC��D|,���|[�2�T�#G�BE眖X���8�Ջ0������?�w:����q�֨���x��û=��[7D����[�S`A�m�.��ށW��W򤹹o�ѫu*)���M���K��I�hz�2>����opBDC*��W�PK�͵���n�/��7|�&d6�@-f��k��N��oڨ#A�"�<!��"� ��?�T����a8 �s�`A��|1��~gY tuvd[����#��������b1�t�;�3l���UY�\M�J���~ƳY#S}��<cY��m�FH���vrL��|�����V�K���,�Yl-�qo�!����}���"D�|)s8��l��)��w�t��aS<ԙd�3��D
�#U��e�|���&V�ݮ�����>�3�odψ��#!at'Ӂ;�~N��w-Qe�b%.)����-o��ļ���h������ �.���;M�E�p%#�s�o����:&�w������ȹ�K���aye0(p̢3}ݤ�؃V�\��9�Q���Ø����+�~����ɕJ1�3�/���J����FE�9��½r�ԛ$}���Nz?a�ط��+"��~��V�#�p	�6q�D�L���WՏ��yn*Ĺ`ȍUR��9>���N�`&��&��%�!J�ӡ��:�?��������/\��3S�<8.��Es��>�&vYX&`L�fE;���4J��� x>͛-=���jE$Ek�G0@il�R�ǣ$((��q���
{a:>ɪ�ỗ{���ܞ���f*����_z;���2l�p��X��͖Q�����~�S�މ~�*D�q��e�~�d*�#�i������ p���%)�Ѣ���U���X6���P_�m�]����`�L�B6hs֡ZZ�￥}��m
+�AD��w[D�hR^"3�W~�"�������/r�d�v`t}kQSQp3�,^|D��y�%^;�B�e.͡s���ߵȪ+�ny����j�뵫�=��Z2S�l�ƃL���D�NSo�g����}��]B;6�5oU�^�Ꙃ���c (�2cm= ��(@%�bx[ �4���L5ƓѰ�%��*~�|vXD�̫��m��އ�U�P��a���K�|�'�T��Ž�]jX����F/x"``��G�~7��(����^$�i���P�� e�M0�i�&� �1S�-�����7�1����z�D��L���
��Ng��a�#MR�Z����R�0[�ɍ#�'��$b`���m7�g=���x)� p�I�m�b�����6�������ōUr��� L9�0��Hz��#Qh:)dզ�{�l���2�p�S�,D�������1^$]L��o�;d4�����k����z{z��f�8������u�����U��cL<kی��Nы9��8�H{�9c߶�-��JУ4�r�}n-��>������r���Udv.S?W>7;8nY��'q[5f}7Sok�3-��8���6IU��*��I��^����n�F�i�}������X�9ғn�����އ1\�xfT�Gk^��$����?�i(���<���o�E ���o�,¡EL�~�oKȿ��N�u��Mٙ���[��l�>�(�V-��8�#!d�/#���O"�^p��ϝ�c�;>�c�e�����ϭz�l�s�E��ԫ4E�֫�	:H�u�Wٶ�#�^E����r�"�L�Mfz��7�9Xq�Ċ�X|>- �>��da�$�^Zh��d��m�v�ӧ[�rS��/uBOp���c��:1�~쀸�0]h=�ʑ*iF<H�g�	���\G���G�:.䡩��滿��z� ��/��*k
��4��
�TrYyS�@U]���	���5)p�e��r���H�	��"7�y���X:!��~�^�O�L"��h�P���Ҟ�+',hV��0o����!�sژF�*��%Ƚ��A���1�x��<�F�!��@���ǰ�Y�,{Pz�c��,G	�=4�&��5<���Q?V�m��[4�r.�k�_�k��ֶ���,�p��	qh���aa	:����.��T�,l�э�v�g�u�hB���(U#�ehCXWM���.S�w�h�K�M��WV'�S��� _��9��e�M���"��N���b�,�\F��s�5�*��Hn�:�A�eү���p�}&���,��Z^���$�b����<�e��!sZUL��Ԗ�!M�G��=|\Y�9�=��sҶ$ڶ�'�u2[W�:N�؏>�)f�@oķ��# bo�0ʙ7)�Z�	F�@�b�&�ӓ#�yi1�D6<ː���am ah���>�z99�L�~�vJ��,��s�.���<�)����$%����K�G��A�r٭�ySR.�1��D�"�`�C�Y�Bpao>�S=y�`2����/�tt�`L���|��В�m�-.^���\m#��Rυ&�����";:':U�}�H���@�l�X5t,��%{9j��]*��!b�O�O�Ly�� tf@T�d7��V�>>�;D��%e�ȩv��WT�v�M�X,�*,�<Piϣ,�����m�>��4l��0x�/�0%k����u(&"��h'(f�hCV���?iK���}����`,@����E�[�܌5�B��n���quR���P�|3%�wE!|K���L�� >%�;�������"\�;5=�Vb���������뻸�p\::��a�I�$�ߞn��E��Y��<}eH����8{�VE���'%��)��R�	<9���u���KoCUR����ڥQ���"�qn���w}4�@���,�8'fH�6�S!���g�5b�<��z)����C���Q 2M~����@V�F���:�@��,!����%$/�<��}R���¾�3�	�8^ �oj�9�=Jc[�6����@5(���S��1���C�3����]y\ OJ��/JE7���bt3*�&d��5BsQ���5z�z.V��������w�#(3'o@`U���x���[Z>:����'m"3������@8+��0��~ M�A��nZ�v�M���	��r�ke�L+�T]��%~z�@౹�%��p`���]:��������8z���Wd�`J���32�ByI0d�}j�9�V�:����44t�&O_��Q��Q���.-#���C��ͅf2*'&��L��K��ӴB4lB���+o���+F��i'����tP�O�PO�ھ��1E����N�-�?��RV-�0�7���S����P�A�8�9��Q�2�>"�:�	!
�;ZuL�qs�7�b��ZŃ�?�\���H^�5�3������Y�Ur`����r�5�Am}�T_Gx=�@n��2϶Xٔ%�ߟ�� �C��$��lyb�\O�q��O-�P.5���z��)_4 ��1��+���Gx�h�Q�v��Y�pP:cP��ؿ�Ti�r��?^w$Oo� 6���1�|���I��??��7qT��+��?n%�Fc�@�`�ί��b�� �mɺe��
1`�D^��ʴ1�j��|�[����Βx�e]���7I
�����0=Ȅū�q��1�4M(˺�x\�~�zǌ��������,\�%Ï�-��Q���{	�]>}�?$��|�IǑg��(ܸ��Qjkg"_Iӣ��x�hK�iUA	���[�I�n����G���;�	ƣT
Fa@�q���f(3N~M�/��|���~�ި��)�� ~��0q��c��C�z�}Iy[�@���`mg�?��5��ۓ�p� d��e�#�?�݊��J� 燓�ܘr��}0H���>�]��I=ڙx]9{���<�-�ߔ�p�� �������:4���b7�f%��7�u0��GC%K1b�=��̈́3Sip�N��3��ǘ�cpQ��j�F���濥׷ʹ�fP��iz�vP�k3]�,�bV���}��,�q,2*|O���ۼ��:L7������"�C*\�5+��n����/��Wl�}
w� e�r��U��B��$Ro�V��Zk|�w ��.:[��֢�Z�Y;LnB�i�"4ۻI$G"�9��
&�. ����A�)����źv�JTS�������m�����^�M}�q���%؏�Ć�������[������n$��!�"�(����f�7�t��b_�p��!��@�&���N��F-�z��Yl&ddV܋d$���mf�͕�.�_��.�dD��Q�E=BX&�00٭���2����B�F��ܣ�]�Q*�WN�{�ԗ�����f�O���~E�	�*Ǻg���$^��'!q�p��P=�$�ut�`�gb����{ꮴ�;�/��'[L�l쯄+�K�]��(���!{�&��!Xz�O3'�3��D�%��s������Y�i��� �O�&��My���}f����&�_tb5x���x9��r2.�y�!����r�uu�|���� ͉swB+W��������G�e*�r���Ó�j�֔�iF
׆�������E�$�Z�
�.��>LG����cǿ-�f��t���.���g��2�V�����8 ��F�̓�u�!��I�ۋ����x̏j��7Q�g��)�>�M�x	��+r����|� �����l^
h	�FԳ)�(�C�c�%a���,�-���Z*���t������)���7�e��TI�����	���p�^B��M���n�wX��	�3'���go�G&8p#r�)���4wQ�\��_\{���-^�,�Z�����FY�m��co����M�1�8�~���\Ȕ��a�;�~h�T�З`Τд��%r��R�H��<ѱ.��=�5���2{s!���'o�7DPo"3�c["��F����D�I0s�8U��2R4k+��t`Ò�G��hd�'k�(�lY���>\�Z"ڊg�+�s�'�Me�"Kw�S6�R������M���M$�	<%S�	��/ug�uE��ی�O xɋ�I�I�����e��C1�Ť�p-
�)�H��!�5% ��MW�gx�y��!GJ���=2�;�|�	��&�Y������4zBԙ)��z�(|����uQ��m��|ڹ�HO��;e ;���2����	Uf��i8a1&�`�o�k�-��DՃ�囘3y�s���;"z�9&�&�V̜Q����S��.�V;>������m"T�D��-M���[��f�NL��j� va�ɏK�yȡ
��jRk�P�JRޔ��Ml����Q.�<�̃:����c��~��m-���\�,�r.��Yh���)VR^��:<��d���5t�_�ͺ ����~<��bOт�9�J��Wܑ�$�cgp�����������Y���N��ZO�M���J�~R��ą��VM>Y�4�N�
:"����&�z�lV�L*sb�Y\3o����Hg����q�����D���I�Q�}K��,V$�}��	�?�	��A!-_�y�x]~�Y�A�$U�<��G8�Ep��X>^ġ|ף���~e��#�]b �!n�Tf��x�Hrg��y�Fp�E��>�ay~`hP��(�Wq6��Ё6/����\t,��)9��}���.��o�G��F�y�����F)����V�:t�lC�B
��K�1kX#�)dl�Q�0��s�kz�/D4�!���F-�]�t�����l���U�虛Q�wfV���J*�$u�GY�v��K�H�t��fҝ��N�QIY�m?-������xk���<�{�&������ҕ���M�%,*�䄱� ����_1�N��ـ��q�&fT�?�d���/ȡFE�t.�+j�ah.]K�p���,}���a-(	�h��g�l�5q�Yu�>�����N�<w��!�:���K�	��S�|\j�R�ĸ�k@��#��w����s�m
uеl!��1�ҫ	>=Yʫ��ݑ�dq��]l��&@�g�ù��(y� �DO1���@ut
hSnd��b�a�jm��m� ��lZ(o>�>�ڼ��#f�����cy���fvn�.)!>BqV}��p�'QRe��e�����{�[l�M`l�5��f���ʫ ��f������Q��A�\C� $��!�j%��d��l����G�l�{5��պ��b��x<�\��qc�����N(&]1٫�oL�����)F7�"p�� �����56r�M�ؙ����e�[�5��!9X���YF]�()׽�a�>@}��奤�r2֬���''w�ן `�����%�X,o�#!��,ƒ�;G�b�^����pu^-c�&r���SeY�����^�*m���z�)��/�m�t�Ȭ
���Em�����鴌��Z��Va��n�Y(�@�oP`�IU!8��i���uZ|e
����2�b����Hט9�m"\��"���tH���S�F�}f-���?꿡��	���Ϳ1�_t�8�L?ApGYl�O���ʶIIǵ퀿d�N��U~;�ͺY\WR��X�����R�Y�3[!�[Q��)j�9e