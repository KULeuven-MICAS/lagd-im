 GITCRYPT �Gf�6$y��	yA0l/zsQB�t�Rȵ�:+I��>�����0���%�l�݇%��;�9�(��[�Ǩ6�^֫Hy�e$��ď��F\�Yϴ+|���ka]�!��5I����d5���U����:�2/��j�G��C,A�l+�m�1iۏp���	[�k�ަ]��bHm �F�+�;?�eQ���қ�Z�Ĵ.�l��p���� x3t�X���ni����ޱ��(��ҧjwP����
zpYs<�XQ��-[ f�ۀ����%�W8�6��E*v�yO�� UP��3�bk(�Ż$?C!9�$��zi�o,l��S�����^�87���zp����#��eJ�����_
@	l2
��2�ɩ�-7��V��#�!g��Q�!-�������8Y��aŮYW�y\אָ�/�!i[B��d^�=�,��U����	 e��]�Qn�9U�s4Y�(Yc6i+�;W��r�|�T���|а�k�t�ퟙS��t�s7�4�H$�V��<�H��;K�Ӫt�י F7fҿ�k~��Kv �;* 5ϮO�@vJ��5�}��NT���v��+�#u���\��X#n���>��/���B���4�Q�;y�RG�Q�ŮDf�D���<�Άd`Z=�-6��Xȫ�v6�	
���C䷿	��-�U���p!�� �DzŹ�P�Q�'� ��HB����K�c��̌>���%� �����=0����<���I)5�Qxb�?i_y�(�C���I�O������7a_#m��?�:��
�����e�|�)dJR���nZ�=_�ݏ+�d��xOCR��h�;�t�9� d����!:ܠ
�h(/`��N8�mf�.�;�a�8�. r�^�"ߴ�O����&�k���&���h%�Z�����w�+�O+��p��+�=���,��|�M|Sw�g�޵OEf��N�V�f��c�����q���!n�q
ښ
��f�j)�u���P�)�V�5ԁ~³�0%����9�5�IQ��\����I:�|�4Y�\�ܙ
,�9��S�W��J���A�g���nc�H�V���Q�E��vD�؀��{e���.dIf�W�$M� ��<��Hb�E��-���_�e*@��Ʀ��H���i9�a�1�08_� ϟG�_^<'wTȹ�vВBeJ��Bqe�ܐ-~�@a��M��`����u�iz�0é0Ŋ��ea��"���Hz�J��� �9g�FS*%�#��uT+��C��ѿ��������?Ö-�%���lҏ�K�$jd3�?D��Sy�x���6j��P˽�f�ݮ1��Q�e&8׃9�)5�!L���

��ۤ���K���,���tMS�5=�4���C�0��kL5�Y�
���A��, ���Y;M���^:A�Ϛt�x^�q
8h)��"�K�`���l���<��r�e ^�_�o9�D~��>y��ޮ�Ї��ȷ����� N6�.KR&�|������\��\A>�G������y�Dk ٬|ˌ�����[�^:��Z��c��oA���#z
��]A�f����u?E��U!�c�ӌ)���/w�G��hD�l�����Ջl�z���^E�����Y+�<YwL�]���f[�pQ�B�tA�l��+O%'��l�*W��A�d=�×װl�1�(-h���O�n�m���6��<��$��̕�y*�ny�d�D���p�ݎ���!��8u~�S�L{[7��/�� }(�r5�A&�Վ)s	��@65��RޣJ*�g�.�+�vK�U,���\l���m��p�<�Θ���-r#�ma�n��'\���
�<D~і�O�p��}�����
�~k�h�`"7�WW�K(9�Wg�`�c�#ðٟ5���\-9yc���@�~5ZOF���z
�t��l����tʰp�N��6E'Ma��Y����Nc9���A���\3 �yt�SR���A|
�l��
�-�R������z�wT�FyE�L��L�5r�(9�������[�*[�o�sjN�⭞"�T�-nyC|�Ԝ�� �s�",P@^k�.�ȸ�+�T�[4�?�+P��xJy�~μ��Y�f��0c=@���d�v���0&io)�~	�iq@\x&�@�����ňl�^���*�s��e��+���;4��Ί��g���/�^J_Qd�m�d��� މ"q!g�'Ԑ��8��1���X�D
�`Y s�ݓFPڷ,�B���K��c����nW�EZ�,�y�d�	��j~YC�}Wf�7het�X;J�E$k���L�D?r�������Q���#�/�\=���� j���&pu�W�+ ��CӺ'=Ye���Z������3�=�� @Đ��-2 +B��S{4R���0ϔ;e�i�y�<�kw��Xzz�
�Z/������|]��u�/����5���3�@N�Ƙ΍Ag��:AF􇣧U�4���Rj�4r���g�p7Jz�te�&Q�E")�ډ:�K�2?@�&��)�~4������+0V0.�}�Pn,<CK�軲kQ��I|�Q+�p�}��ν|�`�h�34������G�T�O�6��}C��S\�rp|ӹ>i���6��99ւIz8�{n��h�:Jjy�ȍ�X��W�?|��*Z�f��z�w��#S�!T�����%c�#�*X:WD�DzX�:A�M�[q�5X;�@��}y�P�谰��2����*��R!�	��0�?���,�i��Բ �?��=~�Q���J�^����?̩a���'*J��̙���Jr'a@�[x,n�?]�ت�Fd��/
I>�}�̅��T������?��殆�+i��1^T����2��S�d�ԗ�n�Vu��2��Jp@�2J��ŋ[�۶�����B5�Miq������W�XB�Ӥ��^熽�u�AR��PC	X�ՃB�2���˥w�g^y�c�X��O��k�"��ocn��D=�?c|in��S��}<��F��͹��X-���j*u�z�[�6]er�����H��gl����qֆL�����ܧ.,��fu@��F�f��Н�_��p(��q�ƽ���u�9�#�~	�#�����%�?1�af�\�`��6�R�
�#t_pux���Z��v�X�PD�Z2u���֎��s�����b޺y��L%�u�V3+��^|)�Bȫ4�S4#5� 4Y��"��XJ����h�;���}�N�J/{��"�j�Xp>.��A�j`��'S�<����aA��w��GDw������nE9����W�#S�Ną�q՛g�st�EȦ;2W�R^|���%�%5�np����UPs ��į7����I
R����ah��ci��UB|�x{����dW;d�&�L[h��`��?Y���|�oφ��`8	fF�k���ۋ�Z�"�98�̘?RL�pc&G�Zzў��W��[d�ݗ���o���71y����@����l�� �:tI�Q����,JU�����&U}�S��� �"5@��:�	���5(B�-�B��u>��_�Ʋm?���4�r=�Z��8��?jpl��N�����Ƽ* �k#��b��|�Y(�^�z'�y❞�V�<ö{�'$�)�*M��B��h�6�T32�?.M�ylrǑ���:@�j��]&��D���D�]r�i��*�e O�v_�4�K��?�\�֒�(Rq��+�
�����q���3�~}���̋-�a���nN��u`�n��%9W˧QQ��`B�Z�;�f����2���r0�좜Z�#=�m������kf+.�T TG)\[ 
�و3��0���S�)��.�\6W#}W<�8'`2$`9�aF�#j�U�0ҿ�hfö���`�/
�mJ=�9�5��mK������͛v2�c$F�(/sSX��L&��H/�Fȳ��[�� dE��-.p��M\$FD?�>P�P�4��>�;7���m"c)��uG�����7��W�л�ZNJC6�`��/�c��UC�_0��h/J_��>�c���R�<"����.��ZX6�Y�ѯ����o�wɄVhM��VY�n���A-3��� ��fY!�z����@�o7��zW�7��K�cɞu�I)�ݛ���{V�+�'��R�ۗj��4.{�M�6�.�߉�Og����}����ҡ�(bч��cE�5v��(�NnΖ� �g+ĵE���	��,!��Y1�����넀�j�=�U�Lh;��ٖ���GҜ)3�]�QE�j׾�\֊�ntd�0��}3�)~!���Q�R���b0�/�5����Y՟Ka���t*�Px�a���8m���Ðq).�X�Vm9�"�|M���2�n5��"���=����"�O��0���T�ߥ"^2��VK\��?(oڮ1���ܑlv�u����G� ��ЍG�/�'�m�����ҟ)��U(���g�	��uA�{�F�n>�:�G*��0-�گ��^�8�>�����A_~��ð���֭�IU�R�B���N2�C�v�x#.����{�+����CGA�vW�y8-��_��fj.F'�r��$*���!�*����VAd��턨��������j��į�6�3]j�s�<U�7������['ͧ.җZ�����H���t�%�X�\/+5��˙��u��KMc{{V�Ƴ�q��	��i�0>y9fbȺ�2dP�/�Eo������t8Ṗ���;c���'z��W�,�~%N��;�i���y6$r�0R��)m�1X�$B������
�_�91Z�C��%�V2��i0ܑ�z������[�A"�TI�wF������Uz/�a���c�p�=�ȶů� q�1q��x��e!�0��_�?g�Q��EJn|�hh��4e���r�nBRqT&jO{m_�,3�D��W<�8��b?�q�C�8��`�fnn]�]��N!� �݀�p@�a�0�����-�W�
��_��>`�E������P���p�Z��#�e���C�m2��.���CbզÇJE��uA��.rJ\�]  ��+�*�g�hY����x^KY<JΓ�G3R^S�4���Q�RJl�����ف��7A��[���R�[-���j��d�� !�;Qb��5'�`�V��2����d���4�R�:T�_�2JG۬�_Ji��Z��q�!��M�5�س�س�W�Xs#!��z�0�Yɨ�̰�|���n��F�9$�v�U��R�Gz�t�u�L��!��M1�O�B@oS�J�}����IC�X��G�o�>/�x�^9��mS��Q8�, -ޗ#��zGU�ۏ���q(#�|��``Q�6�c�U�6�vG�l�9N�d���(g��5�X��/��.�&��$���l�=�ˏ�@��{�I����wܯ$�l3�cUp�W�O4.j���!*�6���{M/�˗_<w�d
Ƒr�&B��ۻ+$w߈�H�/���ЀN%���u)To�+��9�E��7�\���g�=�/2XE���3�M���i �m�����	 ���|Y��S�&vϵ+g6DhF��<9	�g���8BW��D�m^#��sp��0�oɲ���n	���L���.IB~i�o�Z('Q��8��͵�2���i9u�l1&�k�$�B�J�IţK�z(y�ր�|��p�ϖdL�ݼ)�}K>�AM�M��)�X�������;�Բ�������m@��y���;�!�����~�˥m4�80TCMd��1 �P��z�S��+9�T�ˀ'�V|�p���@��c�5r�"8��3����>42I���=��vB�K���r�6<���Ʃ�̱���W��⋛�����K6���eM1�)������`k����v7��_��a%��7o��:{���m�f�J��h�Aw(F<.g�LI�����0k��U��_a��j���;!�Z(�	!*������
�߆q��&W`�,��T�k?����D*�d⡊��rE�|�O��� �x=�T!
�����/fX�ux���ѴQ�k)�,�ز�l�QY
����ʗ����=��2�v��A/�Kɛp�v4;f�#�����I��<g�WP��z�Vl�l^�; A1Al۬��F��r)̌/��`;K�x��D�k'�(��M���(����-���Ƣ���VT�y.�#~|z^ٶ �E���wǘ�N����k?��m�����ϳ�����7k=8u�PsA<L/T�+:�!2�o���X�ۓP�i$1�s]�M��׈�Mm�c*��p��{�4��sB̸>�c1�Q�نk�iv�tD�*ҝ�X+���aX?��L�;SZ?�Ls�-6�Μ�ߏ-𘲭}pz���Y��?��� J�kS��^A�x�rr�]2z���Xm	N�v]
�0�t2���+��w��L�
2'���Հ��w˒S���PW�]������&����l�k�U�=���j�yuD֜�x����L-�rUa?�̋�rM�6U�M�?��+����p��ZR��[D���3�v��u��7�o�:Ⱔ2j0)�����$�ȳ~��n&�!_�-Ug*���2���Y�5���bm��7���)t�Br��<<}x,k\�%��������4�S�tׁ)����AŘ�4�	��3cMrL��4��rק�Z��F��	�L�|sx`Sk���DkU#k(�9�
@>p�R����R���[��<�ڛ6�o}�$[��r7�Y�年����ǻ>P��J#�����J�d����ϋ	/�Ng^Z��t�*�~��"�D���?=�f ٘E��B)�@�P���Re�oa�}}}.�b�� ����/�*U�.�vl���O���h�xin�d9h�>����v�E���U��,1f�eeo^��ݯi��h� �%��v-� �ܠ���]�+M`�Bn���/�xS�[��)��X'��4Y�:����������Kg}da�8&�4j��%��|��� �=���G
���g|oT�����lh/���	=p�Zz�o'�4-�Ǹ��-g$!��5o�2���	���7�{ٖ�F��=|��խ���#�������2��R����78��Bd� ,��@�n��`q�[zl\O��ER�+���"�w�� �J��sxV�
���y����4le�����A�l�7:4TK2��@w;�p
>08S��r7��;�1;��� ��M4���Cr�]BSq�ݞ_"�#1�{���_*�ʎox�� ��rA�]����3�)����;�"��u~L�wζ9k�P�a9��(\���vk��§�[�:jEۨ�(#��4؜��A��2�Fl�|�<�A%�P��h��)�A��5.���H8�+�H�v�o ����:\<W� Kn��K��4�ws�;[�H�������%��|X�����-VS���UY��E&�Bɺ�����;�a�'��}�A�\Ɏ*;P��A!ϛZ��r���P�w-D�4�Of��O����Ό��R;�$��U>Γ;�����̢��P����)%����~��$��;;�AnW.�F���P_��
$� &�)1 �y�B^,3�^�"���MqeL�L����ѣ�����O"�HOf3,�[�O댼k�le`&�z�e��i�1a��Z
�#�n��a��u��'�j0����!���8o�k����6= ���1�����w��[�F�\-���`���÷��l<�)���1"j��/A\ǩ���ҥ���6=>?o@�Aê�}}>h̔�G�ȩ�����*��?Ni��> ��d�z:������M3�C@�hڙ���䝺E��L�v�/a�̦��N���؝s�m�_D���x���ⴎ���Ϻp�h-`� s�z�&���u���
l�}�uk��ߨX���b�E��o����B�D�����B�>����rv|`���k���~������kU���H�.4�7�ԄT%4+�"��lU����tE!�W�C����|2�Ӡ�#u5A,8���W�v���0]S	d��6dϼ�D�KW�F�>�����x��Y[`ˀ���GYn؀݀ E��l����W�5�(sǏ�4eyr;m_j�.lPs�c�/�A���1��d"f�8��%TP2@{��q{Sتk$����M�h�#�DȪ���F�_cx���М�ȯ��)0�y���m�'���0ѻ���A��B�@u�<���K`I����=ٮ ]�p	ԁp��B��0���Nq�"��w�S�W�����E��Q�m"�b�z��`�	F�<oN~�厽)x��`O�*�`���X4��\D��T�&*��B����Ŋ=1k;��D�^�?sʒ6�V����m�ii�u-u<�:���\s���sA% ��2�3�mM�7��3�	4�JA��ǰ��Cj�o<C��Ĳߍ�u�v�ag?��6pHU���ӂr'���������v :����ܶ�c�2"Z����^�늌�R��Pj���3Y8�uu�G�����.s�*8��s��hvK�Y)n�x��׈�t���.���v�Ԩ��
�*�P#���`�P/�L�s�7�/b���⚙�rG����������ZGU*��Q9��'S2;.�����fvSt�S��Y�o�o�,�w�Z��T�}��o�9!{oҕ�.s��-���}����(<�S�����@�045����5�U��X:Y"ێ�?�$=Jfh?��o����5(*���ř	%�^�(��C3�k	�w/����(7qg�RQl��(
��	��\ʼ��lW���C���A�[TF��0,ch%6�f���j^��i�B�*�'3H���|�1	`��Fd��읢?/�JGl�P~��!�m���:�vVq�)J{�t/����C���v[N�yn[������~���>2��x�6��oW��)����('��pw��
ns(Peb�����vC��2��P��z��>��l�������A1�B�JW�6Z���(����[��+�,�$��̶5]dfЖZf�+h^s�#��!���77׎�B�_��w^�@ ӯ=X3�B��,rP���b�|��1M���@��d�[���}��䧦�?y���s;��PJ��!7�^��LS>4�}��iY�9�̅��u5oqy5<y���ՍbYj�T��PHc@I����l�ֱ3-��O�`�4�Z�w԰���&[pOm�|�ކ�%@Q��B�҃[��-g�\ͥ�!�v��B	v��>.�uQ�P^��&|Q��;)��(��O�C��g�b��s����4E8|.7O0>]�
�C���͠c:���2���R��[�uTJo��8