 GITCRYPT �N�)M�mn�p��.����4oD%�Dk��h`�-Y�E����%m��C�	����y�Y�|R���͸Z}����)7��KmrE+��e�=����?�%�_��x{)��80�&���Uğ��M�g�x>�QҮYK��j"���MI�)e����@`�a��n:��u��Ե|H��fێQJa�F���[� !iT�Q\��8a�� �ߐe��ЀJ}���΢���Er�~G��Ĥ\u�F���n��FH<U���)�#��W�#)��$2D���� �^HR)S��d,�|Q�â�l�2!�p{ İ߂m��fA��]$Hw�� �̷��"K�
K�R����4p��GJ��3
l�w,��uW���P�[�NІ��9j��J���X�p'̖�rXF��d��ۃ.v�(�'S{��:� �ɢ辭�/XЯe�9���}T%ҚAB ������QWN��;���b-8%�y�,��A��2N�E��jK-��G6�hT�9E�r~hև����4^�Z���_�khFw']Ci��!���(�\�/�����Ι�
��E���y�3�w��wg�t��`��t��G��/�r��J�����{!k/@�]΅^QQC�hr�z���3���VNw.���A����?�4��	d�y�hN�z���d���O<��k/�8!+ˑjY5�L��ĝh������BQ��m���E��f!���X?_|���,�"&�*;Ĝ�i�i���]�(7��L$���̥��6���b���s������v�]?�Ut���Ք���];��`�vЩd-{��M�`�#[��;t*���r,�!�jb�^l�zA��5�6���#�R���lѮ	x-8%�B 9�=�y$׀I���B)��9�?�ma�_��F�p������389)���`�|�����a���('�]�%�z��2�+O�!���K)�(`��:t����Lav���h->��SF� `{3���{`j抺��L�mh�e*�le�6k�.�	-j�u�[�M�*��*�ƧJI���ܬ���|�DB_�?�&�
ˢ��3�NVl�c;˸ڄ��8N���q�Iq�_L�w�>�	���G��Mĩ3c������"����Y��s�bD���ޑ����&ƭzf�����&��@k�5/�e	�O��g�5aӎ]�y�D]Z�e�� *���3��|y��Ƭ�[{�Fw)�;JU�:e�����S/���@�en�;W_0�"�E;Q��xZr/�~|�-���Ǫ4j���e܄=I���2I9�p�M}��+#<<��lǛ/�
;��s�̣�㞅!h�%���0`ʄ9Wщ�
Ѷ8��u}R��?��x�M��b�>����Eb��<7��\o��2L��X
�M�Tu>j����gDr�������U��_�5�?��_�VƣX1� �F@CS�����Fȹ{�VO��W��!�'0�O"#��Vo�o
(a��S�~�?��8��!X�i�Nq����G�v�P[��?�_n�Q/���H�+Z˛��p�	���O=-�y���׵�]`�o�ZmLa���3<�} 'x�p�}��)ղ[�z�`�����:����΁�<�JVb� �r<upO�_�`�$s�h�	��Ε�+4W+�v�R��z���\UHd����i۰)�H��	b9��Э�����\���33��x�� t�Q%��~@��U�6��ҥ]����%(!`ع�f�=��TXyG����
ӏ=�D�D���N�3c |�WJr�s��(��v-�9�7�ڧ��'U�P!P����R>9fD��yl	��7�]�#9Ջ�ީ� F����;��^����/�_�XqǓ��>�CF�i/�%�L���r7���."sDQ`��)�d���)�\�*�m/bp���p�Se�5-�+� �āL���ۓ
2���c�ʉ��B��]�5Cd
+��v���Ǯ���K{�b�x���4(/d�l^�sʧ�b�v���N�F?Iy�/=����y���j�U+�á�9�}�m�ؤ;��?�O2��~���->a���I�#f�?7ry�w��&|*Yo{�X�o��l�������"�{3my���m�O�E�����!$j���@��8$��t� 3��j��|����E,.��:��<�:	��5�^;�D@���\������g�䕇���##���7x��90���kr���GÌ�&5��ã�����K�����m)�"T�ڋ�h:��Q�@?%u�����o�F��t�R蕵�<���*YD/�9��kD��+��rJ>O��FnV�ZS���Q�xc��P)m3̣���E��G��;V��P�pW��k_�-'�MZ��g����z�Z{�[p�U^�K��}������?�$!;�$2F�b��ڭr���q�v5��3=�٤�Ջ>�/��878������'��#����ȝ��i���2�@�@iK��H?1�4y��0|�w�!�X<z?���Ins֙���5�P)����7YLj���?�
�>�.U�r݀K�n�.D ��8$~�KHJ;��@Mm�s�5=�+�/v�1�c4Q6���|�K̰y�4�6���^��ɇ�چ j�~�?W�(����g��^W���']�U�ᄎ�Y��V�V�mHZ}f����!�g������f �O��IGkb�G&t �0�j(���I䙟7l�a$�q���=���]L��` �z�x�3'p_I ,�eu'>&�ˎ���� 2�@�)hX��L��iP�5�t�Ʒ�7��B���
sf�.x�ɳ�;U�
E��l��T�N3@�`B��*wq�G�/�.pL.��VPE)N:��]ԋY��9駳l^�)#!d�8��`��d�`:���t�qP\�t��'"y���e�?�}�� �T��c�hG��-�i�����Km�J���1.���~� (Bh�r�E��'l�f����u������$���=5{�i�>z[C{#�옚'ٰ����V���ʿ$v*�!^��0��p��p��?x�������w����-��
���0��ywi��i�}�f.�
Y��Z�yjq��l�M��GR8k���f(@��Sgk\�T'].�i�7�,&� BO�1�>F������Ύ��;���!C�T����L�b�t�|�1�L��.�W�L0n����3�L�*��Ɣ����/\���˄�,naW�*%�w$gW���:���?��*��������OEk�t�#�{�}�e{m��:Ҵ��Պ�u�B���c?�����O��k� ��Ŧ?܆,傏��y�����j�"�9n�Q3 >�F�0��E�N�*�O
T�6	A�w�t2�[{�C�4���A�P|����)iCl�Ymy�^��2<����9��Y*8N��C}jY���( 0U�?���![N��!@�|������B��m�㴈���U�2֢'s$�n�la1&��>5�u�Y:�Ί������9����՜��$_�T�{��P�`u��Щ�����չ}�C�0C��iodL�Fj!0��/�8�e��X	=	�t⯙
ӟ�m����i��L;u1��ҷ"j*_���L����#JarO�^���ߜ�g�5�Ř�ڼTty� <%�<���� y,���\�]��ϥ����	f�/��DC��yI�9�v¼4�R�m�t~���vqh}�k	����J�̸硿d����7�.�1�R���E2�����^��@�m7sd����/*��Hz��Ը���a�DE���{�,�uZGv���P���r!Z�<�
)��<�T$VR��߂$ڠ4��C6�:�<�L�6�ޭ�g4}�>Aw[�_�V��zV
}�c�t���I�uE]>}�U^>���Su��č��D	�7����+��
�jf��dn�����C�j�ggױ�-4��_u�<��'���}��/�X�rI��IV�.��S@�E�eST��[��Q[ԽY��uT1HdD���3⋛����44��� ӲȾ���a��5)�����	��AR�N-�y��y�:Mppv������kg�a�_RӤX17Xą����X�����e��آ���\���9@e�rυ�������W�٩�N�{3����αxA�W�%0�V�xq�R��ߑz8��$�=-v�Hs�lB(�I[���Y.��	�B��1s���v�����]Ru�|��R�@�\w�kR{��,X�r>�mm���X�,�C�2���sִ"蝫� ��n�s�S��Õ��I�]�wZ���x�c3�ɤ?�<r~���, &hG<�n�Ѥ9�+���#e� �7+v]�VP>��UlB��S,s\����1q���|p+o�G���	Ɂq�DH~vN��� �+�U>��{-��d��_u�}+�p�M ��� ��T�o~H�(��� ����&nr�C�r���A�yʰ��g��a�Rjw���3�lM?� �b�2�Wa��A��#hCf�\;�����Jd��G%b��d�[i(�-�w��z8�����1�������c����Z��ń�����E��_��Jb|���^�+qJ��5R��y�y=~AõJM���L��!UF�&<�^�dH"	��^:&����K����y��H���،����7���}�l�O��֝�~X����1�~���m��9�G"�n��C2kx�¤���r'k��C�Ҧ"�H������-��j��aj�s+�"H6��}&��%��ٲ��9�T.�,�������������8D�� [� N��r^��3T�T��}g�U�����<ܨ��_K������������?�y�e5'J;t��p��syI�
�q��S�U�޵l�?H�b�5:K:���izd2��l�p��(�-���U�_��o9�UQ�i�6�W�z-4��t���?�t�,��n�)� ,�#c���/�A�y�L'�P:t״�����>Q��eB�~���2A���Ye��ξο&+��g`�B��}�1��ҥ�,^�e��8�����d����H�k�dWA���i* vJ*bO>���*?� P��Ȳ(�,m���O�{Xˏ�y�/'��>���HaI�c[xOn5��(�8,���g�X3A��y79��R�
��.p�g�( j�r ����ˆ�=�	G���>�gZh`��������P�L��-C����r��~��e8��cJ��F|j���"�z�'^�+	��ci���,����%��**���){J�}D��	DNſ���'�)ǫ�#�jNo4E\ċ��>p̥���u��ֆ�� ��nMT��e��T�P�3� �4���fk��;)��2?S[O�#�d����M�
�y��<
�fg=N�`�G��Z�����B=1<�9��^2�f5��f���������t&܌�~Br�=������R�i<���îb?6p�a<�y�����/��uc����"��07�;X$dt|}���v_���{�l�9dNv��z��!F���_�>tMu|h �Dz_�7��	����>����	��C���r�/a�x$j���/$�!gU5��88��M���`-��M������O�y@l���Gd�I���2	l����-sO��f��-m������O<)
�?��_(��jbH�(K��6G��"����d�⠆.��s�4���w�����^�{M�*<o����2Y�,$������ɿi"-�%��x�m������3xj��(z��S6k���u@:d���a�iOs˒k#�nȥ��"���X~�jt�H�Z�e��z���M�t�'�l��Kn��a�4���t�V��+d���+����� �)a,%�b��=l*�C.`���Z���D� �aK5n �¾�ީ@�C�Z��|�.~>$��>Y��?�T�[�k���|N��6D
e��!A,ԮAp̸����f�����/H'�2��u#�u��
E�;Z���6q"$��B� �uK�Y�Q��.cq�Yȱa}�D��U����Q��Y�QGM�ˆ-�P�X G�E�g,"��x)�UP�r5���䚠����Ȗ�ДSrղ
���do����z���w�{����w|��AB��Z�.P�3n�l.�4�mr�0xX� q=0�c�-tB�$�,1�Z���h��%�z:�Z;8���b[�I$>�Ra�,�{[^fH�9�-�-��z���J�}����~N�8*�=��6U;�� �xk���2@�$��#y��]�U���{��>�@��K��/��NMfNqއ�����b|	�:����L��]��8/ۭ/ȡ�$����n!�!S�F�HtYJ�q �Fαw���9��Ф#��~��`�f��� T_�T�+�����Y���U��:у3E��:�ִ	h�C��2O�"��}�
U�j��ԨQ!�$�01�]����#����Mw
�f�^���6���;i9��d հ����P���M\Gt�Vj���B��L?�������z�QI��:.PS�������}qΡA���.Y����&���Ɯ�G�>W��4PRQ�w�G� z4p�����NP���X�k�r�o�=�*���$c�]��E:�>�׿h�&6���95jGP)�^�g��6�	]�.Τ��m�K��1�I�31���!X�[�����jb��w�W(`*�B�9�%%A`��P
�L�y'��I��J|���%�ˏ�}��6]�ͼW�!������1�_e�sa�&����-����Y�z͟e�DG1�c�b_�Q7�7���v��� �.[U���eӍ�yoS�{D"�����c�(@d�����:D�SGA�H&{���?����'�O�֢�@dK�&��<�`ҟ
n���j�z\k倸�1=���Z�2"9Xxʠ�x����c�ER+]��q��9��8����t���a�B��-AQ"�E,U���uM��F���!E���@Ea�إ(*̂��O�a�6NR_����-V�z�JJJ��,\x�C��?���T6f�
p�84����d4)b�O���c�֨b�Ls��,����Ij	� ym�خ����ؖ���0���GLH�><�}ZWsG��Nɉ�ӵ�>��^�9A���Z`�T�Rl$'k�~���}��������9�t��� ��H�9/s[zK
��=zk��c�-��ref���}߿ҏ+�07�"�fG�fF�ͤ�g,��O@�|�,��/�댪�a<��_?�0�Ɲ�K����!�}F����6W����f�W��!�W�UTX�����3�?��aw�N���K����/`
��X�5w*ϝ4��N�yMI��uM/����;�@�ٯ ���'b�� `�Im��hsC[7�Q�W22�/,	e��[b�6��Dij,�M 