 GITCRYPT ֨A������4
�-������H��KꯌP���G��'�O\�wW(E6�����yǟ���[Y��\�B�'wA|�7�${kGЂ��%�D6���3dS+����w������O�
�K�s�M�資ʘ��ށQs9����zX�d��Acr���w����~���k��X��F���U�r�H���l�u&�ɎOR���-Pv���.鈽y,C%�ǃʠ�tU.�E��UBEW�#h�D�\�	[�C�)p/aZ����-�Y�b�l���"��8<%w�Q��?�<0�KȽQY�Ҳjj?;��=�O=�F�Ƀ7��C)�+��˺��ŽX2�M��*��y�ymưt
���-}�Q@G�1u'�`�[	_��_�r�9�H��0,�0GE:�a���L����S��Q!��"O���izP��I�X9q�&�B�u�	*O�Emo!�+ ��:�P��w�w(\� !���jﻼ �	���}�[{e%�������Ω8>60X�����1�#�� =(�E���l�����tQ]�2y�5���ݺ��&����i{�ax��H�Tݤ+�+�A&��U@K�>��f��.7|�o��|�x��2�c������Ĉ~rM�D3)�F*�w�<�FF g��㑫nJ��0�ZO��|�z�:�����nm���h�Tʹ��y�c��<��,Y/� ��Cm����YH�G�~1�-��]80��W�q�˳��Ɵ�S�&�K��Ӽ0	x!��Z8Q��B@�QM�Rz�/�q����u�%4.�l���˔��t{\�>TŻ^�^$�+��1[�+��0:S�7����whK%�C%E�0�	<0�[F>����h;G|؍��.���O�!�f^�{u���@����b�S*��oE�M�a���e������s����4�aU߼f@r�����	QY�Qz<�q_���yo��Q�]�F��B���h�Ȱ�!L���D�	kX%ع��)y�}���e�(WX�j��
�h�y���Ft�����ਇQF]f��._�-(�`-����(Q�I�׷٤���p�j�Ģ�X)>��cI~�ma9ΙF綰d�5���g��բ|ج	ɏ������TS,4�!��#��ʬ�܄}7.#�\����=LVvg��+J
L��%���i1�"�~��E~HO#VQ"U����1��9���g��A��mB@s6�|�3O#��a��&�,�Y�c�&j�fN<9=��ѷ�g"�*�Wi���%/C��v�̤9�����͆����YUǳ����N���������w���䒜�<����jB��O�2 �է钀���J��9����T:-.�#l���M��4�? �6�������@@u�AQ8}�P1Կ�-�+���e7���OV��|
dV��C��K�U�l��s�<U!�&/�r>�ɾ�4�x*�`iZP8��N�q�f��w"�(�j�R�O�)�@a��*=����s�l"���}��(ť\��n�:_��א�(� �(��~y�,0XE ��5s�V3�t���-	���3����J�V�z�7L]�մ~�QXK-P��DfkA8���=Ů�0à�T �<
3�׈��0N�����0�뗑_*/�۷C���%��{Uޢ���ᜥK�Ƥ�P1�k����̿���F�"��:2j��6"��c2ةSE�0B(�FV�Qf`���,g�g2؊�+����۩Xɂ��]c4{}�����KA+��a!��^���	H#c��f��j*R������?D::��!����N��[�� �$u�˕���z��N�b��ʙE�nE�P8�符!��D��gvS�A��֘"�]���H�b�3���Y�����jH=mE�\pv�����O@MAo��bi��2C,����ˮ��P���l��$��q�+θ�O�l6D�b�1����P���Ţ�,.v'�}�A� ;&��G�+�''B�C���_I$�\�E��:�r�ݒͳ�V� ���غ�=�x��q*�6p��F���Nj�b�[��ؖ���Ci&�wt	ueV�2wa�c���₣A8e�gt��~B��F,Ӣ���XR%g�;�y��!q�q'��7��
܏�*ѻ<��1�]�{�����@���>+1���?clc�J�t�/]�9�T��'@^#��}�臝7�f� �7����! �!ʆ:�١Z�x��	��-��*�hkڬ'��$a�ox�+zt�4`~+*�� ۃTm�>��1�($�L�~n�!��']G�ºl�%��TVկ$��Ji�^�"���<E��E|\���i��;P��R���v������Y�N�1�Ym�����������ײ=��&��n����_��YL0<�����}�eT�Rvu�������/&���h&]^�V~)��2Ϛ��~w#�����t������[_���*+���RF��4pRN��--S�#��p�Y�9!;<9���?�F\4���[�� �q��q�&�fJ��� ���r���^/si2�6�6�U[�x'��܏m	��l6+��v#�ʭ�r�^"P��$}G�3�oh?�Y��$����`�5�D=d�s�8�WkJ�|��禷fh<�����\���Y���WɒT0r�)IԽ�A���5�3g\t�D�^V[���Ji ��%����9\�ӷ�c�)�kưy��<-lӱ��|�`*�.eܜ�0�NFD�1+��{it���MǴ�������u> ����`U��Ꮌu앟�W8�XP��A�O���Α�!�S��*`
��Kd`�-��œ�H�\w��$!���Zf�u�JT��S	���'�+��3�4rК�R����:�3�"t�_+�N�(���wi�ղ�m�w�K�r�IQ�xGϬ�j��F�U���;B� V���s�X�}��ܝ����i>+}���"��܂,�o�H�6�g����ךi�3b�}B������|�f���y iM�x������.�}�{?��e����rl��|ؤ�LO�b">�RG^�V6:�"w��\7�3C&���)����*	��� ����Ս�Z�y�p��k�Z9#S03�ޙiB�<=z)��+2� �ľ5i�����wv&�Ǣ��QSg8�:cBmcu~�;��@3oĪ?��oQ7R6�b
F�T�g\u"WQm�����HY��.�_��SV_�%�1�˗���>���i�FX#�c�-�#	�e��c���.T" )񒄀����w=��/��$2���a�4D<ln��X��-�N���Pt���/��r�ͷf���pw�฾�/�L�ͅ N��1y?1Y�����S���ܗc&�-�}�g8�Mh�\OfZe�\<���&R?�2�n`4�&��ݼ���>2����U�g���m%�ف�&��U���
��{9�%���
cC�?��~��+՚jP����x�"k�E^����t��nc�Zy�����)�.�P�'4�Zdj�v��C��0�{;���@�*(,ʮ��(5���i�
V�!S_��[yD�7[�t���E��n����ǒn���by�Is�
�1YG]��'��f���	���`��G����r/>D���V�6Gk�Y>�E��
x�iD��lhG�W��K�6QR�d5h�dOP����x�V�a�AV��<�i*P䤇I8
�A��b�C?Bi�R� }����&?W�g
�t<$}Y�`�'�1�mWQR����~ב��
�����8Xfő�ן�=�V����R㛋�L�j�I���e&���%BM��l���+�*1���g����窒/E�P/~WV�[���*r��ُzKb؆V0?DS������`�;A�ϝu�a��p�zc�lB��pq�Fr�;u��ĦG��5����G;����,@��֬��q�4�!bA c��)0Y[}�������.��VI�`�jm{%J�	F4N;}כ��敹���0�/�rT�M݀P��|kv��1��*}[f->r�lI�/"�`�?����K��$��`u˅[��ʠ�����,��e�,(�}ޙ���ܝu��S+5˹Fd��+�,J3g,���_�AJ�DPMR�~����D�xɩ�I��>2Zi��{��Y"}�Cr~��6a���jc*����k&]����G�Dl@_��5*JL���䡮�ML�Z�h�+R���r?S��_�=�>l���Az<��n�<<j�*9-`γ�P5�w�;"`��+Ѓ\U�z���}���e�o�Eo7֋�C��l���?����^x�`J��4�����E��&�-��>��K�������G��m��5���ne����h?5��y��ybԉ��e;��y��.�Wt�U)X��;v�r�-�SNX��>��r7ԨF3�H�fГA�6R?pB��A��;��H��]c��=��������ۿ��3љDH'�Q_���9�K�j�C���(��9�f������t��M#$k,�[;E��a���e����C��N1�.����i�^�	�Ke�n��V�3�Xb�Үl0�}j��LL����V�񄫒j%�A�0��&%|j�Bd�PLŪ��
�Ċ�8��{$O���U��a�j��i�.; P)�쵕>��� k�i�����5�E<�R�v�Kŀ�����|u�qna�g�<z!1��+,x�M��e.��ۏV�Wġ7�B��Jͩg��M�!g��:rVp�w�-���j�^��ؼ)���b��C~5�O��O�*����4iw��"�9��ŇΫ\�&w������_+T��q��� �����[��˷��*�"�D�\2�v1�Rp���ʣQH6�]1�<�b ����W��oYƵ�	��N���r���)�3;������e���^qX=�b�0O��&�-��,U~N��l��ݬ1��0!��2��@Ҥ
�z�H��_3ϸDF��C<�.��lK�u�4��$�*�.���b�� ��b}���HT7��+Z?K��Q��g]��B��.P����uaad���
�r�b!gTTf��C�+0P h|�����R�"�>�9'^��o�*�Ǩ�"}<`,�\(�R5�$ I�����xO�H82d���k�{�I��@T��~���� {#7חA/�OG(��U�{�o~��0���h8�,F���w��S{�+7�>	w�-ܣ^KޝO]�8�ޑ�SL��-�m��a�Y����R�rQ�bl,`i'�𱜫,�.׏�%�D]%xt�6�}�v#�9A�ܶ�8��8�b@�h���[�#^El/9���Dt�Yv�
��<oep4�A�Miuu�/��$�Lj�9�٥a�Ҋ�ʘ��9��{&��$�����`q�K��=A��]v`����뀡����4?�����u�e>��K�g^à�:�%�z��M�l�
,+G�����OQ��V�I��'�c;	��<��#x��V�� @ݓf*���o�M��,�>,6ǀ8_-iH�Q�ܷp�g�.gͯ�#��ħ��K���
<�U72�,���_���k�K�#ֺM��RW �c���,�e�6#�=�
r���혠��F|a�:0��SAj��9���rymS�?Y����*soc�֪���p�K���)%�c��Y�@h,(��T}.?���ɯ�~��E��~�� �_*Дܢ<���Ad[L2����#z<FaZ�RA�>u��|�����A�Fo.�*'��'��G$��RҦā���ݽ;�����#֏�(��o����VpQV��&d��n(x����qf҉�2~Ja���p<��kEEJa���ܴ�.�ե�a�{.�<�����Be,vPx{����:�N j
���6�im6Te���/a�Gq¶�cSiY���6$�i��3=�-�\� �����=�i�v�$`��Rv."Q���C��� t�<z����ޤ���DG�L���#�i�Y�t&_��|#70��S:�*��E�O8K���xu�Sغ��m/:��5��ߍ�t��ݫ��+�`�}�j�|���G>�K��c�`Qfw��` ����~ǡ�����E�|���?d��~���R[�~��+��1��b��םby��ަ�Iy��"�M�o�j�@�-�l�^2�cd"�#���0��o[�X��x�p6WG$=Ls�(R)RI��p�
V�Q��(�r��ܦD�%}��L�<3��K�����,% ;�|ߌW���l�]a�Mܨ�x�(怟�x�Q��6�h���0X�H21T.r�s��5p�I	�?\�i:��>��x���CDi��.!Ʃ���\�T̈@oK��KEB>�޵�y���WJJ3�͎�#����^fIQ+�����d%�{�'5O�J�P�M��s���&S-�D6Ajꡰh���M��f����Xs�k�Tt5�'ae���3^��ͮp�Z�u�>�#F�����}u��YM�L�!\wߐ����搸:�{8�q�i4g��M��%�l�_�X"��G*�*���у���or{	�I�Ԡ��f������-�q��\�8��:�4i�"0��B祉�5B�i�1 �6�����%v�I�ҹ��c�S�b�Աv�{�v������(�P���������>��4��
ЭL���<�W��S�ʷ�>,�R fv%�i��ʊk��rMCv�ej���p[w쌓n��".*�m���$��� ���\�V��Q���`��m�U�IkG���h��/ဘpPĝrbP�M*���W �,�����!� �7�Z4�ǃ4��(b� n�*���X�����o� Z<���={;�I��,�@ۣ ��&����Dc�q�_xS��{7L�`��Y���G� u���z�A_ͻ�Q�~�i�@%��z�jZ��o�<���M��i�BP��i,߻�)�Y�����L5%yJ�H�YG��"M³o�&T�M@�9����x�+�cב,��tJ�r��p��#xl}��6I~�|V��e�\�4��|��*%���($�h~-����L��9�ʫ�tɬ�ߓ-����25��<9���V�*�rkV�&����`.*�~��'#���o�Է�a%@�]-���|nS�S�}v�jO��ǀ^ H�}���4Ϯʈak�P: �4>�6֦UtR7.�NF`V�,=6+�v�u=M��o�u��6�<�쩨yn�+0#V��n\�9@����
�Kͱ���{��Ѯ#/�L8���F��9;��
�U��t�P*0W���biZy�κ� �U����h+}�Tn����N��#qz	�l�#���Zݯ��B��>O&�l�O�ɔ�j۱$C��Ɏ��cF3��~���L�	iV%��������K��O�Y��vb��x'���]79�)��0&nss�g�`x("���g���g��w $���lH�ש