 GITCRYPT �No����+�6nn��{7y�lQ���讕bK�U��w�z"eS��~���K���{�!qE;����T��v"�;��w���aS�0�}�]��U�-�b2>�HIG��dz�+���<D��l@8��r)=�N�a��� D� b�{-0(?�h=��$�Jئc��. �0ɫ��?���zM���0Qv��k������I��c��������	d�mBZ���� �#Y�z���_����,V�Ko�×	K������8��J�5�!�l��c����K�3L�o�(^}@���ȃ�,�^�4ۡD:�D�J���7�xQ��{(o��q�����	ا����N���B�j�b�=4ږ/�,�ނQ����u&�w�cv����/~�i(Uu�6Q��o��S�E�Axad��*�*�F��e�!���t�'�Ω:��=�j;0D�1Z�����ӯ1B����#kv`��Z�P�y��~?���?�>?�O [���㡂���a���f�&��?� {絣n�%ǰA(z����$5l�R�D��E�E۾	�:� 8�_x��FĚx\1�C�������Y�HܱF]�|	^�oBX�L\':7M��^\��>�I�����.(:&��ņD�/"��nΰZ3�ͳe��CP���5~p-қS��:����2�{h���Toz1z�7p�:�F|y�J^9�!y�;�����(=�H�3se�������Y�4�b5J3��|)�q�P��L�8Kq����x��\\�{�_���(=R�cމ�dءp�&?*�A��&���p��0@�眛=�yy�CׇŎ�5�\R�I��ƚ��{�#�+%��	����G:�g��t�����^��1�A8!��.7G��l���]���=\��g�*h�	s7/ƨ�t/p����hY���K	�t�ޤݻO�&�4m5�R��"X�`���15��������SF��&~��|�@�͑���6�V�\	�����/�]��U:�\�^��mq��D�L�^�w�$,���>6DJ#
1=����ܾA�6[
C[��U���F��
��n����!�+T���F��=�x�{�l-`��������fNF0��BY��mn��қQ���kqkK���hij�f���U������9��LuOm��PuH��Zc�K"pI�_���u?��j)<@��xP\qD?�����'�<	��6E9[^�AMO^b��h��V�������P%�-���LQ�Y���y�7�G>��\>j2�����Ѥ��n�����$��ͯ������NrN��ѩ��N���j�@J2�*A�2�=�xĄm�ǙPp^�F��;�:�L��aþ�iu��c��SYC_TK�D`��W?��6�4��A!\��?xB�?Udx�����#s`�B����ۯ#�����C������TD��G�`Ϣ���ܒG5�v}���r	-L���gu�4��&\����# �-�MI�#<Z摮�ۇ_��q�D�9`��tȚK����_��^����|iۇ�ׂ��wb���8����ᣏ��i���w��=����"IYN�
O�ۉ0�����4i�7~���.J���ԟ'�eF�Ul�A���4?�h���C�Q%�PF�$�9.-�+�a8=��9�3�N�U�1+�$��X~Z0��Un��4����7���)ڬt������o"P���^��b<��FQ�Qx����$�GЉ�Y�@�p���M��kϱ
M���eB��4xp���\:�7�D�<^�]nغU7��h^_yt�Ik
H����/r����+J~��ِ{D�'���n�\g�?FBgާ�;����_��M� �+?\�_�NAie[-t	-��,���f�W����7v}����(W�ꡨwUP��4���3��j��"G�4�/�5�_ۓѻ�܁���{�,t�Z���(YZ�8�����8K�]���>qP#�h��x�RC�e�&	�Һ� E��yML�*�q�B�T�@V��$�!3�O!$ '���Ъ�$��7�!�w*�����a�Х�-y�ߠ���s1���}�#!j�4zHq!^��u��D��-�hm�Jɾ���"�A��e��=c\OP�5��+�,���/�7��P���T�1'M.��S�1��u�]�4��Ј�.g�_[<�:���m���0Tj齨E*m~�كά��ў��D_9�w�e���a�9�n�<봢b1Z����wՋV3Hn�YRM�`��n�
P��_J��oK����wz��%�S_F�4�.'{bT۪���&�Ul��:�c	H1�g�� ��'����Hhz��!6�sP���e��7�+�zP؏فJJ�HlW�7G�y�Ň��"�E�����z��ĠO{䜚~r"�y���q�0�^o����C�~����O�Rc�#�F1�_E,L�ds���fY�=�w�W,r�؀��1�X�>�+sݴ ����v���� g��Թi��8曂~��83��RWX,��iW����9Fʩ�yZ���P9���O`��k�问ԉ��F:J䰬���D��,P���6=A�a�'����F�(�=2�p�=D�Q0=3:���������^�n��H�c룲���w,1�E��u��W�~ևEʨ�pܽ���)T��o�1
�Y�� <s�CԘS8���m)�j���ά��v�k�%g@[���o$܁�����*E7��>;Ȕ.�����:*P5�l�\]��HQ���$���h����Mb�sY̕�ᲆdg�>�$���[�H,�����i�}3��`"�'�j�AZ��6�����jS���zc���ͮ.XYY#9<U��P�3�RmL���p\�d��:��x��q_ӳ��V'� "
�W�������>�hߙRɘo�r�_��%����n^r�Xyz+^>ח��s�+'���3	3_�k�
ܾ%�w\��~mdP����~/*�Ì
�`H&���\���'�-�}$=^e'��Gs�g^(R+>R �}�T'9H����4�x\W�*f�ﮃeژ���o /N'�Y;�P�:����mج�f�U눡h����J�� @7�nfP�,i��Zj^{����Wb0Ű(�deĨ;��6������Y�`l��5�ְ$��~*����D"�3���,Xiܕ����&M%�xS���1dKl����6��UM�-�L`�K��7�I�['�S���L�
�_��h��ZW��x���[��I`����6�Xl��)��(�ԆC��.uu;�d��1�����Po��Ca�&*�nb�+JB\��p�lZ��[Q�C3�{N�dH�+�Vq2�\��ݕ����Nk��r>�R�?A��D��AB778�OO\Y��[n�Mh�}����8:��R���=]jP�k�o-���R��s����8�p���X����H,�/:��߻�?Yr15�Mq#,d�7�����(���^��}���Ukh<����)+r7!�lcFA�\��q��7iP]�N*�=Q�F���Fn�u��Y�Ϧ�?�vX��߸�}���,9��'u�`6;e�������~\/�����2˲L�Y1����ڕ�=���Э�	0�TR+�;�v4���	:2#��Kӆf�mE⢆"��נ��/�xE�s�Gn�r��lr���"�ƥ��f�FE<Z(�)��/�E��Ӎ➑	� f�CA�l7��.$?;��!D��:�sHt��[�h�r�D��-���N��P�@�|���e�x���aT0���'�����@��T�@�[(E��0�I&w��0tbU�N��a�!�m���e�6 �t�pQrY�^���t�Ȳ�mn��]p�T�"�
��B�	j�y��t�%E����݅�X��p���Q{'� �dN���Q<܈�\n�Ϡ�d- 7���B�@�,N �(>�_��k���~m��E��Є�8L��	��6~qp��Ƚ�\4��m�|T6��h��B��׮Y���gd���:ǽ�Ycq+�qU�$��L%Lr�M"/y�Vp�P�{��"JT�G�d'2�&x*��ާ�lBQZ�<�=0�_w1�e��&E����Y�i��U�c�?����Y��r�mdPx*�E�b��Ml��es�.��9��q�0�)��:����	U�	M$�w���-W%��FԩB��:<�DY5z�d��MP{��vnI�i�%�/C�\�ʌ�C&������\��5=��}5�}�V��WV�=O+0���9n�O�zm��[!�?M ��̉�WO�D�.���<9�*D �d�V%���]5��N�q �����4mn�c��
\�&�Fcm��r��6�t���K`!��9z8r��ˤ��a0'��D��a�'�pM�ȴ���4����=�<��&����7�r@cS�Y#s��*b���߶�K���j�Wɀ]B��
�*�N���w��bA�Y$)�2�;�P���:l#� ��L��S^ %(��)$!��𚙨���R<��b�%��bH���k~�C7]���f���� �8X����B��qy}4��{�Ԗ*�������"��V+����\	5BB��S�^�f`���e�6��(����mY#�`%��G@���O"F صI��s��cn�]�m.���*7s�g�>P �,H��\�3�i�I�R7�-�d���I�3	��vE]�㮢������Ir5G��i{1�ڹ3L����q�,�˶B�CPr��2��"H&�g�ޒ��oJ��s����{�b���B�'ۅ0թ����+g&�zB�.��u��k��i��	V�	��榢���#�H��l {0�'�)Cs���)V�㯾�#�� @�<2EY�	�Cv1���O�5'�>�g�k�vµT�s񪼺��J1.5뵂���{�N�ȇu�Av���lX�:XD�BA�f-(��/�`�0�t&��Fy�~A]��=�Ҩ��Փ�4a��A�FN`�!�jT���G��fQC^.�5�������� ,d�}C��NT�\��S��~���,e�������#�jݜSih�_&�d�t��mN���Z�s�2k����%�r���0�'��Zk��\N�>��L���tH��z}'Ǚֿd����4[�{l%�*��aN$��!���K��	)����੕څ��؛������ΘƁi_v��>YR4x6#=�?,,VƜ�O��`��S����2�c��_�z��5hXf�ݣ�1z*���
�������X���Pr�2��;�B�U�Q���q���=��} ��\(z�y� ��>��fY̢�%��(�/q��a)��f�z�,�\�؇j106LI�f�e�#'��� n�^j:�*J�C�D2�Myb`,�'u��rq�ړ3`��;�kU�+�<�9�I��l8wHr�A ;��{�fz��LXR�����x�-�H��N���1��Ȣ�^װD�gD�������[5��*�HEܚ��a�c8=@+���e�X:��;�#h|�W��#������ǝ?��� "��{1$H�1�M�����Y4oX�����	�H��:�6`�����j�^���oz�`�.Km�w�RT�H�y��	��|�y�(B��_C[1�t�U@кZ��9ª���g����8E���iRg�nb��GE֋o�2Hk+�@�JS� R�؍��������f�
Ѩ�mS�C�o*Nmq�:�+P,�g'�E*Z���F�G��o��q]
 xV3�ܞ_f8�R�|\��'�Kt�%o�FP�.����q0ݸޖ̿��	i�Oa����n�� ��u�u�GZBc;0o�Y�@��S�>�ͧ��r�v����S�G�x�ݰ�� J��Z��dQ��%�*�  �+�	B^|�a�B6L��G��A<��Y�R��Lw���5˿&~`�c�C���Q��!��6�s^{�ǅ�Pa�09��I�MU!��R>�Q�d��ӆZq;��)nz#���@�K�ď���͊69[A#�E�B�ci��Ŕ=����-Rpop[��|�.ݟS��kь8)�:f�O_v��[��;�`cv�o�LM+��',�p|*7���&�d���P֢�P�Q�����u�eL�3��: ZP�ʫ��p߹�M��C�t	�X�U�Ԕ�l��C�3Ǘ572�x����_
��<P���u��W;�A`�դ��Z�����I��tLLuaU�CV�z �{���PnC�_T���\���� n��ɾ���TY�<��=�d9���wp�5��?�1wl4ڻ^�8-���6<BSs�����#$/�؏۱���T�e]�9����[����=?�ㇳi�	b�J��vբ�z�I�w�3������b�f�����ȱ�����2�A�8ya�M��|�w).ˤ,R�&ӷ�����JJo����`�48(����b< wJe_�|�,���]^e�̇z=��q#�+�Z�ư���S;�/~++�,˷t�K�F�2��J�K}~D���n�7�I��E��Y�.�c���:�`������ c`��l��f�]]3�<R�R�$��!$����0�oH���
�8m�c]�-X�;lD���,�@Ove�O���k,Lg�9׀w��+A��+1����lT0����b��Ml\9���bQe_��.M��e	dsQL���m�x�o�m�}�C�-Ztؾ!�h�?v���R�'�ƭMp	$zJ(ED�4������cZw���%v�L��g�����ؙ��z���S�O#�l�k Y[��Y�i~5� XrP���2;A���%#����?�xD���4\h�<��N���~�E���c����n1��1/�e�܉���N�2, �F6���]^��v����D�_���hv<��Q�	��W^�0��=�����7��t\��|��V,%�c|�3�^Օ�.P^>�4�0M}Ԇ�b-@HF����VZ�,�D�h�Q��1J�:�{a̋�Q��چ
��'����=6�uO��k��;���$Ѳ�dH����zD[�x2_D�Ќއ�T�e��{�"ع)�X��fWi���Մ���D�t7b�5xjo�R��eO�! P�����:�ca,=x
sE�H���Pɪ�#w����fKq�V���#;2��ዜv�m�k����
��8s�	0Spx*5z�gX�l��ׅ� ���'����O�<d�ߋ�R���S���XX��=ڋ��T�4������:��A�Fu�~�L�2~�|aN��ʵu�|q$���s�nmC�\�%��,#c@�)��Б�@�֥;ڶ�h�������R��>s:	fFu+p}Zx>MF�ONĺ+�������W�QXh�_�;�R#�