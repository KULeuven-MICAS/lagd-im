 GITCRYPT V���c�1]K3?J�h�g�+���á]�f����1Y���{����9�K��^�:�C?��Mߝ�
�<8߀*^��/��1(��#&���2�BD���W�	�gtv��I 02���nޚT����w��_��Mz����S�g��hr�.a��)�ivJ��b{��񧸄�(����嶅\��Ou�M��3�7*E��&�¨ïr�?�0$<�G��F[+!Y�lMH0�5���DV֕�$ x9�y!2%���|�����Ϊ���]��Ϟ���4�lJ�_���Xj�'��"qWL��DL��'`�H�&�ˑ?�",T����h�'lCG�r��s�U����^�������m�Q��ď��0�W�˞�;I$kEŁ	D.��߮BM��3�:D�����l}
������k|Ș��ʈ�����:26U�\�ؘ��.s}I���x[��Üazˡ�_�:�?�JO�P�:b9V�#��]T��f����� �= �K1A��������'n�78�מ�J�$r��҄Nu���t T���3iq9S�X���-S���%�R�e1�5��y���V4�aYe6�m���<KY�>��˻��* H�=w��ε�Բ�b�1+5�U���̪ݫMR�0����>>�))�Ǘ^�L͍k�%V�:s�/j�F�B4Q���R���U��Kԃ�n:Y��3�s9��`p��@��;��k���'4(L��%㬈�j����&�l+)��&���x�u�/�����x_�����a�
NfD��d�W�v�̻���GH:����XꄩBu5U\��Pw�;5���7�?DV�|��I#�j; \��<�`K�vZ���XLRH8N���_K�K�q!��fK�c|�2��v���'0� � ���g<A�Fx�YQ��g�w��YY�b�Ŷ����7� +�t�g���?�&u�U���p|�,�ڱ)n,��W
'o��@P5g��{_���Z��h}��+M="u*����h���a����i|�V�<a-�?>��lW�w0D4ăfk���������Ō� ��$\�/�v�G��S�=����6E������p>���\��LqW���D��#�Pv�D���mKm��M��7�z?.�3l�C�T�ߜ�a=�u_�Ӧ�G��e�M=���=��}uL��[6f�[���1�s�o�����S���<0X�^�\�@�;�y�С�q:u�s�+�]wO<F�q,��-��'��ᛧX�J���F�"p���h5;}vj�X��@@�L�d�_��)�P5�I*x� �
*����syx���o�0u�~��	{��Զwl��a�D��i$H
��s2�_���zf��.~V���c�󲔖� �7g̑��}(}9�c�'�i��p��Y��qT���+[��\嗫oḶB淲)"X|CBz��Z�t�o�NFlh������9']�q��^F��x]��d���N�����v��4���=Zl��|�m����=�~��9(�=y���Mw���$�{��k��pNI��.��'�O�k�0;>t�E+Rf~U!쯢�\�.�ʢ��+��̓
�dK�������_5�hn��y�u�R;Hw�mк��G
�F���GK���Y7�h2���|BJ�Rn"�˹$F�m���Mk�8D�W�\j��O���]H�r����uBe�%���4WQ!���`�K�zKP�DU:�rDN�ZB�Ȋz�*��-!L�l�Dt��	h���ߓ��ĩ'�:s�����OB�+�\FS�D�n`����*on�p�_ȡQ�{�;"Fʜ�)6&1On�J�`=��VA��3J��l��1)�����u7��!���u�����۞���#tm�q͡��#F k��rE���&�	_iȻn��1Bt��#59���O+5���5/UQxig�-{���u2�1�E|7ŵ7�_���y �t��`#�+S�&�/9I��I��������9����Ә;�w�����
����z�,��t6��&I#�u&k��u�I���f]����>�G{Jn����56!~y�_�S.d��mq>���82\ޱ��\(�:�k�R�\�^�}����n�
1$9ݳ�KDݟ���!��w����!n���D�b���A\I��y�M ���\���3�6@ܑ�H����\UҢssǼ��gR��rC<����EGe����ґ�Y�t0d�Ԓͦpʰ���)}�M��mjf�5����`ʏ�bV�ΈYr�	h=a�=@6��J&���yC�n�D���KǦ��Ӻa9:�q�=����hw���#��"�l�Dm����d���ߔNK�.Xqb�L��8�,��?�����Ӭ3t�2��r<�5���_{I@�Lc~\8��L��h:�����K�	:&:�jTɨ���b�� ����Nw�D1��X�6���8f�sӦ�{��7�AV10�Ӆ���6�3?|. bh�>ޛL9:���TYKO�(0�E���Sd�p�i��.��[\d2�p[���#����GPv�*��}��O-鏓��������/��>�/w�	��~'5}®��}~�����`1��6WUJȕO���<(�\��b���Y��mh���L�x~���#�'*���wZ�72o#@����Y��Ԩ�%d��miT���,|	���`�O6s�= K�ŬW�
�x7A4혹҄���Y��r&�.�Z��M� p<f��{���哱��dv:;<e�2Ԉ��m���ő�v��R�pUx���jȓ���ޒ�ם���	<9�D-#O���M�����	�YHż�Z~�x�cSʎN�V�Eq�8T�8)va�F�-)�ڟj]��}g:O��׋J�&�Z�8�KV�a�t���5��e>9�������{>ڬ�����<㙰3l�Ж����^����M�`�j('D�֜Q�1'H�H�^�%�$�m�~�=DDQ��m�\��!�XO'�!�J,id2rQj�/��[��\R���ɶ�'8�.>9���AW.�w�Dk\z��#��m�/�)ŃdO���~6QZ�(��?���p>��//_�q�S�'�6���.� o�H�M�����t��[�Mr�J}�t�>��E���8�o?n�TU�v���7���b��[i�kC�G�T_Y,�VC�W9�;���]t��4���������w�e%�u����K��-�M��V��e��ϡ"��C���j\1��ۂ���!�;�&@���7�N����:)P15	�
�7o���js���P�.�/\���GΉ��g.�����=(�)�:I�2HWN��9��^��������r'�J��N�`���|˯���F���k ����r�hRE��΄��I%&��J����V�Qܸp8�Z�2������oOR������&��'M��k4:>�^�xC�
��ex4�@�=�K�߶� (�lT��}��VR��� 2O��zZ}��'������:��Έ�[m��g�w��BS���@��ؠ7��?�!0Q�[�Q��E�s��M�A8�b���������_s�Q�oA���AO1Ɉ�DI����S���q&B��8M��ң��2�C�HM����>҇RCA�]�r�ȯlxs���H/#/fM05ѽ^ã��ĕ�P����ߘ�Ň��4�'xs��(�{��?�z޾y�%[R�C�~��a���n�E�+Χ���"������<0ҏSh�*�=t��/��Xp�^/�0�ǫtCe���3���:�;�R�/����&�cB�v�QQN�lT6'��6�ٶ�#����R�4tl`�
/�6�_A�^Oy��w�x�\8����U����o ��D�b_ȯ�r�fEof�e�ZcE���-[=h���ط҃�/}k�T�;T���aC�^v#w#$Z�K�~�Dp���\~�}H�Y�3�}t��ԋ�gHI���/��;8�McB�v$xI���y%LHx2d��ZY�S������cw�*]y�͕�!w�"�L��3��Z��q]���(VB�+L��"�x�Uc��pY8)=���n JbXp��w��t���fɲ�y6���V����Լ�cB��.�A�p�O¿��µ!�:lb�����)xBk�R(�zM,�OI<��7R1�cD��'>m�nѬ�����WxB�T�F�J?ǧ����1ot������/`���މOX<��[�6!����(Y�#�(�{1�K~���/o�9��J��PE���n�X	��0��U\^���O�!v΍c)�U�U��<V+`QI:���]�~1���������S9+��c�7�7i��}��o�{�|"��ab�!���g����7�l@�Q�e�TH����.x$;����
y7{�|[	�a�܈K�:y�'�8g��c�q����&M�>���X!~�L�j�ɬ��B�P�k�tX�~�̮��cn9�VJ+��#��?|����t�h��4�ٕ0�e��%ru9���R{�4�mGC0h�}�+��hE�BB�L����E�h���7�BS�[��{����5e�֑7��dM����u����|�4�շ&6����1��w<2�Uj���uKk�d�Y*�7����,8�U<gwWV��s����������	jB��E���qV���~���?8�ՌtQ���x��Pн���x�k9�gXG��N���9nɸu�ЙZp����n�~��]�1����[�m���.u���=��E�w�����ѫtz�ND�	:"{N�6�":t��"> ݆�2Ϛտ~'y	���5�w'�r��������#��e�!�����>����#Q�MHE���Fw,�)��p`�
v�D����<�L�SSs��d�x�K�X'�D���?\0BC��5ra���=�bl���c�"�0c���j��-���f#�}+��vݬ~T_$�g݋�LZ�G �;���N���`B�*�)+F���{����3~nY%'H��<OCN�-d���L~:� X�^)Y���!�G��O���M���֥�q��=��
��� {b u4{��`�Ga����=Cp*�`8�b�����tc��dh'��Y^�T�8̆	��!�����<	}&�)�}%I�u���\��1�s�2��LENٿ�09��K�ش�Ovb�]�������[��k$���=�dI�%��g=� ��\۹�ign幑A�8e1*�\V��/͆5°�t����2�:�A����<�p�ζHG��":H� �A�l2�X������9@��!�d2-}G���[���]ѷ�w6���(f�|�8����!0A�-�Ըr]���F]������{b�g~��j�Z�~%2�:�W�!OiKnq��C�>Q���'=k)r����y�]z�@}u#	R��E�\~lC�_�'�V*�* -� ��ٍ���A���3a�RL�_�ш���X���[m4��B�S34ZM�gHt+��E��\+�׆�kq�����L�jj%�]�*�h0�'��T�z��X����Sی��
��L��_���+�7.4���Eٗ/RF��OO^ܥ;`�+���9��ml��c�N�w�x�������o���5��fvΑ�%�I�$�^��j�n��b�p���:�qc�}f$���$�ؤ�BNT!�V\���kܔ��:έ&=�-����#���,���Q�������WL������%4m���C�i��

�K��(��i�<��L��$���Z㦼��P�p.{�1����,,.0��q�~�6�B��48�+ �<�v�m���}^�V�`�n�5�F�� kv�Ӳc�9���Dľ��;g�7�A1��Δ���B���1�Y^m�c7�%��ޓ��{Њ6I��v@fNj y+��ug�PW����s�>�{Da����o�V�vɡ#YHToX��1�_�k�ɅHG�^��.{��Q�X��E�>� �0��W5BVq�c�5qLza�g:0^��v(}��2�ߔ����>��L;�UyR��w��)����� h��qG;���!f��뉈c��
��^���;	;�,Dޝa�֓�CZ�Xb�^����� 2�\4�qM��ۙ$>��9}��<S���)�Q�ī�������pF�1��G�K��p)�ŷwO1gJeg��6��Q���S�f�]�?��P��=��t04g�,5bW�sq.���ܚ`د�l\Od.����9�N�lg�og���v�ҧ�>��F��T6rUZ��uwm	4�����!` �R;��3DH�����é�Ɯl�8����<���Na!Y�Pg�r�K9x�u=`a?/:��~�
P�;�n�x��>����!�
Xb�_z����d2U��r�qk~gh�O��B�Q��
�[0fIOg����XA�|i��
#��X����A�O3��s���@�c� �<�-�JQ'�|���c�-����\\˵�ͪw����
�M5(Jd��ߧ|W�;�7��3�{�e�����⸂F����������SU*=oȕ�B�W�n��(�˶�|�f{g��#��)�7tC2�j��0/� -�iRg��H߫��@�Q+����@5f�/˒�\���Ӏ,�~�������0_�A�ϕٶ3����O\k38��+J���S8�b�o��'p=n}nHly.i�`u>�@*�W� �z7��, t�8�X�*\Ό����Ԯ� ���B��������0d�̹��ʤ�;K�������G��=�R%�ہ��Y�i�'��vC.�����"Q��rK%��b�	���F�ԩ�s�p�)������k"�D��<��\�|��*&���P���0G��&x�>q�o��b��>�@�˔��� {���P���Y,�cC3o�7��V�X��?��l撦KlB�P����~�RE��;��lmC.Hց��X��t�&�:=�/q��ܪX�n�>]�5�}n
|�r듐��nZ�+���0���l�5�G�~b�,Gp^[���ao�ӄ�kH Q�vk�+��ROl���;��bƯC���T��b�? �WD�\d��3�U���C�
B�(�z��c�qwd=��SXs:�E��O��xz:��H �r���Ę���ݗ\F�Z��,h�SDa�����ͭ��]ZS۪��a���R�o!�Ҹ�g��MIEy�s�̈��K4=k~Dq���m�8������=��D�٠/��<a++p4�.n�ˣ.����7<�߾)��.kGI�FװRB10��OE���g^%]��s�u�b�,�9��f�e?)lp`��7�x���Ɔ��R����q�´���]��Ϭ}]�w���1���6��!7���TLⰹ�Jk�n�*�y��Q[�